// ---------------------------
// Nome: Jorge Luis dos Santos Leal
//	Matricula: 417466 - Exercicio04 - Guia06
// --------------------------- 
`include "clock.v"
 
module pulse ( signal, clock ); 
input clock; 
output signal; 
reg signal; 

always @ ( clock ) begin 
signal = 1'b1; 
#24 signal = 1'b0; 
#24 signal = 1'b1; 
#24 signal = 1'b0; 
end 

endmodule // pulse 

module Exemplo0044; 
wire clock; 
clock clk ( clock ); 
reg p; 
wire p1; 
pulse pulse1 ( p1, clock ); 

initial begin 
p = 1'b0; 
end 

initial begin 
$display("Exercicio 04 - Jorge Luis - Matricula: 417466");
$dumpfile ( "Exemplo0044.vcd" );
$display("Tempo - Clock - Pulso");
$monitor($time,,clock,,p1,,p); 
$dumpvars ( 1, clock, p1, p); 
 
#376 $finish; 
end 
endmodule // Exemplo0044 

/*
TESTE				

    Exercicio 04 - Jorge Luis - Matricula: 417466
    Tempo - Clock - Pulso
	
                       0 0 1 0
                      12 1 1 0
                      24 0 0 0
                      36 1 0 0
                      48 0 1 0
                      60 1 1 1
                      72 0 1 1
                      84 1 1 1
                      96 0 0 1
                     108 1 0 1
                     120 0 1 1
                     132 1 1 1
                     144 0 1 1
                     156 1 1 1
                     168 0 0 1
                     180 1 0 0
                     192 0 1 0
                     204 1 1 0
                     216 0 1 0
                     228 1 1 0
                     240 0 0 0
                     252 1 0 0
                     264 0 1 0
                     276 1 1 0
                     288 0 1 0
                     300 1 1 0
                     312 0 0 0
                     324 1 0 0
                     336 0 1 0
                     348 1 1 0
                     360 0 1 1
                     372 1 1 1
                     384 0 0 1
                     396 1 0 1
                     408 0 1 1
                     420 1 1 1
                     432 0 1 1
                     444 1 1 1
                     456 0 0 1
                     468 1 0 1
                     480 0 1 1
                     492 1 1 1
                     504 0 1 1
                     516 1 1 1
                     528 0 0 1
                     540 1 0 1
                     552 0 1 1
                     564 1 1 1
                     576 0 1 1
                     588 1 1 1
                     600 0 0 0
                     612 1 0 0
                     624 0 1 0
                     636 1 1 0
                     648 0 1 0
                     660 1 1 0
                     672 0 0 0
                     684 1 0 0
                     696 0 1 0
                     708 1 1 0
                     720 0 1 0
                     732 1 1 0
                     744 0 0 0
                     756 1 0 0
                     768 0 1 0
                     780 1 1 0
                     792 0 1 0
                     804 1 1 0
                     816 0 0 0
                     828 1 0 0
                     840 0 1 0
                     852 1 1 0
                     864 0 1 0
                     876 1 1 0
                     888 0 0 0
                     900 1 0 1
                     912 0 1 1
                     924 1 1 1
                     936 0 1 1
                     948 1 1 1
                     960 0 0 1
                     972 1 0 1
                     984 0 1 1
                     996 1 1 1
                    1008 0 1 1
                    1020 1 1 1
                    1032 0 0 1
                    1044 1 0 1
                    1056 0 1 1
                    1068 1 1 1
                    1080 0 1 1
                    1092 1 1 1
                    1104 0 0 1
                    1116 1 0 1
                    1128 0 1 1
                    1140 1 1 1
                    1152 0 1 1
                    1164 1 1 1
                    1176 0 0 1
                    1188 1 0 1
                    1200 0 1 1
                    1212 1 1 1
                    1224 0 1 1
                    1236 1 1 1
                    1248 0 0 1
                    1260 1 0 0
                    1272 0 1 0
                    1284 1 1 0
                    1296 0 1 0
                    1308 1 1 0
                    1320 0 0 0
                    1332 1 0 0
                    1344 0 1 0
                    1356 1 1 0
                    1368 0 1 0
                    1380 1 1 0
                    1392 0 0 0
                    1404 1 0 0
                    1416 0 1 0
                    1428 1 1 0
                    1440 0 1 0
                    1452 1 1 0
                    1464 0 0 0
                    1476 1 0 0
                    1488 0 1 0
                    1500 1 1 0
                    1512 0 1 0
                    1524 1 1 0
                    1536 0 0 0
                    1548 1 0 0
                    1560 0 1 0
                    1572 1 1 0
                    1584 0 1 0
                    1596 1 1 0
                    1608 0 0 0
                    1620 1 0 0
                    1632 0 1 0
*/