//ARQ1 - Eduardo Botelho de Andrade - Guia03

module rand (output [3:0] s,
             input  [3:0] a,
             input  [3:0] b);

 and and1 (s[0],a[0],b[0]);
 and and2 (s[1],a[1],b[1]);
 and and3 (s[2],a[2],b[2]);
 and and4 (s[3],a[3],b[3]);

endmodule 

module ror (output [3:0] s,
            input [3:0] a,
            input [3:0] b);
            
 or or1 (s[0],a[0],b[0]);
 or or2 (s[1],a[1],b[1]);
 or or3 (s[2],a[2],b[2]);
 or or4 (s[3],a[3],b[3]);

endmodule

module rnot (output [3:0] s,
             input [3:0] a);
             
 assign s = ~a;

endmodule

module f4 (output [3:0] s,
           input [3:0] chave, //definida apenas por 0000 ou 0001
           input [3:0] a,
           input [3:0] b);

 wire [3:0] w1;
 wire [3:0] w2;
 wire [3:0] w3;
 wire [3:0] w4;
 wire [3:0] w5;

 rand and1 (w1,a,b);
 ror or1 (w2,a,b);
 rnot not1 (w3,chave);
 rand and2 (w4,w1,chave);
 rand and3 (w5,w2,w3);
 ror or2 (s,w4,w5);

endmodule

module test_f4;
       reg  [3:0] x;
       reg  [3:0] y;
       reg  [3:0] chave;
       wire [3:0] z;

       f4 modulo (z,chave,x,y);


   initial begin
      $display("Eduardo Botelho de Andrade - 427395");
      $display("Test LU's module");
      $display("Chave: 0 = OR / 1 = AND");
      $monitor("x = %b , y = %b , s = %b     - chave = %b ",x,y,z,chave);

      #1 x = 4'b0000; y = 4'b0000; chave = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;

      #1 x = 4'b0001;
      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;

      #1 x = 4'b0010;
      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;

      #1 x = 4'b0011;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;

      #1 x = 4'b0100;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;

      #1 x = 4'b0101;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;

      #1 x = 4'b0110;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;

      #1 x = 4'b0111;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;

      #1 x = 4'b1000;  chave = 4'b0001;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;
      
      #1 x = 4'b1001;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;
      
      #1 x = 4'b1010;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;
      
      #1 x = 4'b1011;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;
      
      #1 x = 4'b1100;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;

      #1 x=4'b1101;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;

      #1 x=4'b1110;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;

      #1 x=4'b1111;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;

   end

endmodule // test_f4
