// Exemplo0011 - BASE
// Nome: Vitor Angelo Lima
// Matricula: 451621

module test_base_01;
	reg [2:0] a;
	reg [3:0] b;
	reg [4:0] c;
	reg [4:0] d;
	initial begin
		$display("Exemplo0011 - Vitor Angelo Lima - 451621");
		$display("Test number system");
		a= 5;
		b= 10;
		c= 15;
		d= 20;
		$display("\nPositive value");
		$display("a = %d = %3b", a, a);
		$display("b = %d = %4b", a, a);
		$display("c = %d = %5b", a, a);
		$display("b = %d = %4b", b, b);
		$display("c = %d = %5b", c, c);
		$display("d = %d = %5b", d, d);
		$display("d = %d = %5o", d, d);
		$display("d = %d = %5h", d, d);
	end
endmodule

