//------------------------------------------------------
//--- Avalia��o 01 - Nome: Jorge Luis dos Santos Leal
//--- Matricula; 417466
//------------------------------------------------------
/*
	  0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010 1011 1100 1101 1110 1111
S0 =   0	  1    1    1     0	  0    1    1    0    0    0    1    0    0    0    0	
S1 =	 1	  0    0    0     0	  1    0    0    0    0    1    0    0    0    0    1	
s2 =	 0	  0    0    0     1	  0    0    0    1    1    0    1    1    1    1    0		

  ---e) Montar a equa��o simplificada do sinal S1 pelo mapa de Veitch-Karnaugh:
  ---- (~a~b~c~d) + (~ab~cd) + (a~bc~d) + (abcd)

*/
 module saidaS1Mapa(s1,a,b,c,d);
	input a,b,c,d;
	output s1;

   assign s1 = (~a&~b&~c&~d)|(~a&b&~c&d)|(a&~b&c&~d)|(a&b&c&d);
 
   endmodule//saida s1

  module Teste;

	reg a,b,c,d;
	wire s1;

	saidaS1Mapa saida (s1,a,b,c,d);

	initial begin
	a=0; b=0; c=0; d=0;
	end

	initial begin

	#1 $display(" Jorge Luis dos Santos Leal ");
	#1 $display("letra e)");
	#1 $display(" a | b | c | d | s1 ");
	$monitor(" %b | %b | %b | %b |  %b ", a,b,c,d,s1);
		   
    #1  a=0; b=0; c=0; d=1;
    #1  a=0; b=0; c=1; d=0; 
    #1  a=0; b=0; c=1; d=1; 
    #1  a=0; b=1; c=0; d=0; 
    #1  a=0; b=1; c=0; d=1; 
    #1  a=0; b=1; c=1; d=0; 
    #1  a=0; b=1; c=1; d=1; 
    #1  a=1; b=0; c=0; d=0; 
    #1  a=1; b=0; c=0; d=1;
    #1  a=1; b=0; c=1; d=0;
    #1  a=1; b=0; c=1; d=1;
    #1  a=1; b=1; c=0; d=0;
    #1  a=1; b=1; c=0; d=1;
    #1  a=1; b=1; c=1; d=0;
    #1  a=1; b=1; c=1; d=1; 

	end	
   endmodule//teste

