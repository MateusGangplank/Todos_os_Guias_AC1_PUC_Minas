// ------------------------------------
// Guia 05_03 - 3 bits Multiplier
// Nome: Alyson Deives
// Matricula: 416589
// ------------------------------------

// ------------------------------------
// -- 3 bits multiplier
// ------------------------------------

module three_bits_multiplier(s,a,b);
output [5:0] s;
input [2:0] a;
input [2:0] b;
wire [3:0] c;
wire [3:0] d;
wire [3:0] e;
wire [3:0] f;
wire [4:0] g;
wire [4:0] h;

and AND1 (s[0],a[0],b[0]);
and AND2 (c[0],a[1],b[0]);
and AND3 (c[1],a[2],b[0]);
and AND4 (d[0],a[0],b[1]);
and AND5 (d[1],a[1],b[1]);
and AND6 (d[2],a[2],b[1]);
and AND7 (f[1],a[0],b[2]);
and AND8 (f[2],a[1],b[2]);
and AND9 (f[3],a[2],b[2]);

assign c[2] = 0;
assign c[3] = 0;
assign d[0] = d0;
assign d[3] = 0;
assign f[0] = 0;

four_bits_fulladder_nor FBFA1 (g,c,d);

assign e[0] = g[0];
assign e[1] = g[1];
assign e[2] = g[2];
assign e[3] = g[3];

four_bits_fulladder_nor FBFA2 (h,e,f);

assign s[1] = h[0];
assign s[2] = h[1];
assign s[3] = h[2];
assign s[4] = h[3];
assign s[5] = h[4];

endmodule //three_bits_multiplier

// ------------------------------------
// -- 4 bits full adder with NOR gate
// ------------------------------------

module four_bits_fulladder_nor (c,a,b);
output [4:0] c;
input [3:0] a;
input [3:0] b;


halfadder_nor HA1 (c[0],carry1,a[0],b[0]);
fulladder_nor FA1 (c[1],carry2,a[1],b[1],carry1);
fulladder_nor FA2 (c[2],carry3,a[2],b[2],carry2);
fulladder_nor FA3 (c[3],c[4],a[3],b[3],carry3);

endmodule // 4_bits_full_adder_nor


// -------------------------------
// -- full adder with NOR gate
// -------------------------------

module fulladder_nor (c0,c1,r,s,t);
output c0,c1;
input r,s,t;
wire carry1,carry2,cout;

halfadder_nor HA1 (cout,carry1,r,s);
halfadder_nor HA2 (c0,carry2,cout,t);
or_nor OR1 (c1,carry1,carry2);

endmodule // full_adder

// -------------------------------
// -- half adder with NOR gate
// -------------------------------

module halfadder_nor (s0, s1, a, b);
 output s0,s1;
 input  a, b;
 
  xor_nor XOR1 (s0,a,b);
  and_nor AND1 (s1,a,b);

endmodule // halfadder_nor

// ---------------------
// -- xor with NOR gate
// ---------------------

module xor_nor (s, a, b);
 output s;
 input  a, b;
 wire temp1,temp2,temp3,temp4,temp5,temp6;
 
  nor NOR1 (temp1,b,b);
  nor NOR2 (temp2,a,a);
  nor NOR3 (temp3,a,temp1);
  nor NOR4 (temp4,b,temp2);
  nor NOR5 (temp5, temp3, temp4); 
  nor NOR6 (s, temp5, temp5); 
  
endmodule // xor_nor


// ---------------------
// -- and with NOR gate
// ---------------------

module and_nor (s, a, b);
 output s;
 input  a, b;
 wire temp1,temp2;
 
  nor NOR1 (temp1,a,a);
  nor NOR2 (temp2,b,b);
  nor NOR3 (s, temp1,temp2);

endmodule // and_nor

// ---------------------
// -- or with NOR gate
// ---------------------

module or_nor (s, a, b);
 output s;
 input  a, b;
 wire temp1;
 
  nor NOR1 (temp1,a,b);
  nor NOR2 (s,temp1,temp1);
  
endmodule // or_nor


// ----------------------------------
// -- test three_bits_multiplier
// ----------------------------------

module test;
 reg [2:0]  a;
 reg [2:0]  b;
 wire [5:0] c;
 integer i,j;
          
// instancia
 three_bits_multiplier TBM1 (c,a,b);
 
initial begin:start
      a=0; b=0;
 end
 
 
 // parte principal
 initial begin:main
      $display("Guia 05_03 - Alyson Deives - 416589");
      $display("MULTIPLICADOR de 3 bits\n");
		$display("\n   A   x   B  =   S  \n");
		$monitor("  %b%b%b x %b%b%b = %b%b%b%b%b%b", a[2],a[1],a[0],b[2],b[1],b[0],c[5],c[4],c[3],c[2],c[1],c[0]); 
  for(i=0;i<=15;i=i+1) 
  	begin
	
  		for(j=0;j<=15;j=j+1) 
  			begin
			#1 a = i;b=j;
								 			 
  		end	
  end 
end    

endmodule // test three_bits_multiplier

	// -----------------------------
	// -- TESTE
	// -----------------------------
	//-- Guia 05_03 - Alyson Deives - 416589
	//-- MULTIPLICADOR de 3 bits
    
    // --  A   x   B  =   S  
    
    // --  000 x 000 = 000000
    // --  000 x 001 = 000000
    // --  000 x 010 = 000000
    // --  000 x 011 = 000000
    // --  000 x 100 = 000000
    // --  000 x 101 = 000000
    // --  000 x 110 = 000000
    // --  000 x 111 = 000000
    // --  000 x 000 = 000000
    // --  000 x 001 = 000000
    // --  000 x 010 = 000000
    // --  000 x 011 = 000000
    // --  000 x 100 = 000000
    // --  000 x 101 = 000000
    // --  000 x 110 = 000000
    // --  000 x 111 = 000000
    // --  001 x 000 = 000000
    // --  001 x 001 = 000001
    // --  001 x 010 = 000010
    // --  001 x 011 = 000011
    // --  001 x 100 = 000100
    // --  001 x 101 = 000101
    // --  001 x 110 = 000110
    // --  001 x 111 = 000111
    // --  001 x 000 = 000000
    // --  001 x 001 = 000001
    // --  001 x 010 = 000010
    // --  001 x 011 = 000011
    // --  001 x 100 = 000100
    // --  001 x 101 = 000101
    // --  001 x 110 = 000110
    // --  001 x 111 = 000111
    // --  010 x 000 = 000000
    // --  010 x 001 = 000010
    // --  010 x 010 = 000100
    // --  010 x 011 = 000110
    // --  010 x 100 = 001000
    // --  010 x 101 = 001010
    // --  010 x 110 = 001100
    // --  010 x 111 = 001110
    // --  010 x 000 = 000000
    // --  010 x 001 = 000010
    // --  010 x 010 = 000100
    // --  010 x 011 = 000110
    // --  010 x 100 = 001000
    // --  010 x 101 = 001010
    // --  010 x 110 = 001100
    // --  010 x 111 = 001110
    // --  011 x 000 = 000000
    // --  011 x 001 = 000011
    // --  011 x 010 = 000110
    // --  011 x 011 = 001001
    // --  011 x 100 = 001100
    // --  011 x 101 = 001111
    // --  011 x 110 = 010010
    // --  011 x 111 = 010101
    // --  011 x 000 = 000000
    // --  011 x 001 = 000011
    // --  011 x 010 = 000110
    // --  011 x 011 = 001001
    // --  011 x 100 = 001100
    // --  011 x 101 = 001111
    // --  011 x 110 = 010010
    // --  011 x 111 = 010101
    // --  100 x 000 = 000000
    // --  100 x 001 = 000100
    // --  100 x 010 = 001000
    // --  100 x 011 = 001100
    // --  100 x 100 = 010000
    // --  100 x 101 = 010100
    // --  100 x 110 = 011000
    // --  100 x 111 = 011100
    // --  100 x 000 = 000000
    // --  100 x 001 = 000100
    // --  100 x 010 = 001000
    // --  100 x 011 = 001100
    // --  100 x 100 = 010000
    // --  100 x 101 = 010100
    // --  100 x 110 = 011000
    // --  100 x 111 = 011100
    // --  101 x 000 = 000000
    // --  101 x 001 = 000101
    // --  101 x 010 = 001010
    // --  101 x 011 = 001111
    // --  101 x 100 = 010100
    // --  101 x 101 = 011001
    // --  101 x 110 = 011110
    // --  101 x 111 = 100011
    // --  101 x 000 = 000000
    // --  101 x 001 = 000101
    // --  101 x 010 = 001010
    // --  101 x 011 = 001111
    // --  101 x 100 = 010100
    // --  101 x 101 = 011001
    // --  101 x 110 = 011110
    // --  101 x 111 = 100011
    // --  110 x 000 = 000000
    // --  110 x 001 = 000110
    // --  110 x 010 = 001100
    // --  110 x 011 = 010010
    // --  110 x 100 = 011000
    // --  110 x 101 = 011110
    // --  110 x 110 = 100100
    // --  110 x 111 = 101010
    // --  110 x 000 = 000000
    // --  110 x 001 = 000110
    // --  110 x 010 = 001100
    // --  110 x 011 = 010010
    // --  110 x 100 = 011000
    // --  110 x 101 = 011110
    // --  110 x 110 = 100100
    // --  110 x 111 = 101010
    // --  111 x 000 = 000000
    // --  111 x 001 = 000111
    // --  111 x 010 = 001110
    // --  111 x 011 = 010101
    // --  111 x 100 = 011100
    // --  111 x 101 = 100011
    // --  111 x 110 = 101010
    // --  111 x 111 = 110001
    // --  111 x 000 = 000000
    // --  111 x 001 = 000111
    // --  111 x 010 = 001110
    // --  111 x 011 = 010101
    // --  111 x 100 = 011100
    // --  111 x 101 = 100011
    // --  111 x 110 = 101010
    // --  111 x 111 = 110001
    // --  000 x 000 = 000000
    // --  000 x 001 = 000000
    // --  000 x 010 = 000000
    // --  000 x 011 = 000000
    // --  000 x 100 = 000000
    // --  000 x 101 = 000000
    // --  000 x 110 = 000000
    // --  000 x 111 = 000000
    // --  000 x 000 = 000000
    // --  000 x 001 = 000000
    // --  000 x 010 = 000000
    // --  000 x 011 = 000000
    // --  000 x 100 = 000000
    // --  000 x 101 = 000000
    // --  000 x 110 = 000000
    // --  000 x 111 = 000000
    // --  001 x 000 = 000000
    // --  001 x 001 = 000001
    // --  001 x 010 = 000010
    // --  001 x 011 = 000011
    // --  001 x 100 = 000100
    // --  001 x 101 = 000101
    // --  001 x 110 = 000110
    // --  001 x 111 = 000111
    // --  001 x 000 = 000000
    // --  001 x 001 = 000001
    // --  001 x 010 = 000010
    // --  001 x 011 = 000011
    // --  001 x 100 = 000100
    // --  001 x 101 = 000101
    // --  001 x 110 = 000110
    // --  001 x 111 = 000111
    // --  010 x 000 = 000000
    // --  010 x 001 = 000010
    // --  010 x 010 = 000100
    // --  010 x 011 = 000110
    // --  010 x 100 = 001000
    // --  010 x 101 = 001010
    // --  010 x 110 = 001100
    // --  010 x 111 = 001110
    // --  010 x 000 = 000000
    // --  010 x 001 = 000010
    // --  010 x 010 = 000100
    // --  010 x 011 = 000110
    // --  010 x 100 = 001000
    // --  010 x 101 = 001010
    // --  010 x 110 = 001100
    // --  010 x 111 = 001110
    // --  011 x 000 = 000000
    // --  011 x 001 = 000011
    // --  011 x 010 = 000110
    // --  011 x 011 = 001001
    // --  011 x 100 = 001100
    // --  011 x 101 = 001111
    // --  011 x 110 = 010010
    // --  011 x 111 = 010101
    // --  011 x 000 = 000000
    // --  011 x 001 = 000011
    // --  011 x 010 = 000110
    // --  011 x 011 = 001001
    // --  011 x 100 = 001100
    // --  011 x 101 = 001111
    // --  011 x 110 = 010010
    // --  011 x 111 = 010101
    // --  100 x 000 = 000000
    // --  100 x 001 = 000100
    // --  100 x 010 = 001000
    // --  100 x 011 = 001100
    // --  100 x 100 = 010000
    // --  100 x 101 = 010100
    // --  100 x 110 = 011000
    // --  100 x 111 = 011100
    // --  100 x 000 = 000000
    // --  100 x 001 = 000100
    // --  100 x 010 = 001000
    // --  100 x 011 = 001100
    // --  100 x 100 = 010000
    // --  100 x 101 = 010100
    // --  100 x 110 = 011000
    // --  100 x 111 = 011100
    // --  101 x 000 = 000000
    // --  101 x 001 = 000101
    // --  101 x 010 = 001010
    // --  101 x 011 = 001111
    // --  101 x 100 = 010100
    // --  101 x 101 = 011001
    // --  101 x 110 = 011110
    // --  101 x 111 = 100011
    // --  101 x 000 = 000000
    // --  101 x 001 = 000101
    // --  101 x 010 = 001010
    // --  101 x 011 = 001111
    // --  101 x 100 = 010100
    // --  101 x 101 = 011001
    // --  101 x 110 = 011110
    // --  101 x 111 = 100011
    // --  110 x 000 = 000000
    // --  110 x 001 = 000110
    // --  110 x 010 = 001100
    // --  110 x 011 = 010010
    // --  110 x 100 = 011000
    // --  110 x 101 = 011110
    // --  110 x 110 = 100100
    // --  110 x 111 = 101010
    // --  110 x 000 = 000000
    // --  110 x 001 = 000110
    // --  110 x 010 = 001100
    // --  110 x 011 = 010010
    // --  110 x 100 = 011000
    // --  110 x 101 = 011110
    // --  110 x 110 = 100100
    // --  110 x 111 = 101010
    // --  111 x 000 = 000000
    // --  111 x 001 = 000111
    // --  111 x 010 = 001110
    // --  111 x 011 = 010101
    // --  111 x 100 = 011100
    // --  111 x 101 = 100011
    // --  111 x 110 = 101010
    // --  111 x 111 = 110001
    // --  111 x 000 = 000000
    // --  111 x 001 = 000111
    // --  111 x 010 = 001110
    // --  111 x 011 = 010101
    // --  111 x 100 = 011100
    // --  111 x 101 = 100011
    // --  111 x 110 = 101010
    // --  111 x 111 = 110001
