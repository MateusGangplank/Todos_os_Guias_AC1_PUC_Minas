module Exercicio01(cout, s, a, b);
	output[3:0] s;
	output cout;
	input[3:0] a, b;
	wire t1, t2, t3;

	meiaSoma HALFADDER1(t1, s[0], a[0], b[0]);
	somaCompleta FULLADDER1(t2, s[1], t1, a[1], b[1]);
	somaCompleta FULLADDER2(t3, s[2], t2, a[2], b[2]);
	somaCompleta FULLADDER3(cout, s[3], t3, a[3], b[3]);
endmodule

module somaCompleta(cout, s, cin, a, b);
	output cout, s;
	input cin, a, b;
	wire t1, t2, t3;
	meiaSoma HALFADDER1(t2, t1, a, b);
	meiaSoma HALFADDER2(t3, s, t1, cin);
	or OR1(cout, t3, t2);
endmodule

module meiaSoma(cout, s, a, b);
	output cout, s;
	input a, b;
	xor XOR1(s, a, b);
	and AND1(cout, a, b);
endmodule

module testeExercicio01;
	reg[3:0] a, b;
	wire[3:0] s;
	wire cout;
	integer i, j, linha;
	
	Exercicio01 FULLADDER4BITS(cout, s, a, b);

	initial begin
		a = 0;
		b = 0;
		linha = -1;
	end

	initial begin
		$display("Exercicio 01 - Douglas Borges - 417889");
		$display("Circuito Somador Completo de 4 Bits\n");

		#1 $display("       a   +   b  = C Soma");

		for(i = 0; i < 16; i = i + 1)begin
			a = i;
			for(j = 0; j < 16; j = j + 1)begin
				#1 b = j; linha = linha + 1;
				#1 $display("  %3d %4b + %4b = %b %4b", linha, a, b, cout, s);
			end
		end
	end

/*
Exercicio 01 - Douglas Borges - 417889
Circuito Somador Completo de 4 Bits

       a   +   b  = C Soma
    0 0000 + 0000 = 0 0000
    1 0000 + 0001 = 0 0001
    2 0000 + 0010 = 0 0010
    3 0000 + 0011 = 0 0011
    4 0000 + 0100 = 0 0100
    5 0000 + 0101 = 0 0101
    6 0000 + 0110 = 0 0110
    7 0000 + 0111 = 0 0111
    8 0000 + 1000 = 0 1000
    9 0000 + 1001 = 0 1001
   10 0000 + 1010 = 0 1010
   11 0000 + 1011 = 0 1011
   12 0000 + 1100 = 0 1100
   13 0000 + 1101 = 0 1101
   14 0000 + 1110 = 0 1110
   15 0000 + 1111 = 0 1111
   16 0001 + 0000 = 0 0001
   17 0001 + 0001 = 0 0010
   18 0001 + 0010 = 0 0011
   19 0001 + 0011 = 0 0100
   20 0001 + 0100 = 0 0101
   21 0001 + 0101 = 0 0110
   22 0001 + 0110 = 0 0111
   23 0001 + 0111 = 0 1000
   24 0001 + 1000 = 0 1001
   25 0001 + 1001 = 0 1010
   26 0001 + 1010 = 0 1011
   27 0001 + 1011 = 0 1100
   28 0001 + 1100 = 0 1101
   29 0001 + 1101 = 0 1110
   30 0001 + 1110 = 0 1111
   31 0001 + 1111 = 1 0000
   32 0010 + 0000 = 0 0010
   33 0010 + 0001 = 0 0011
   34 0010 + 0010 = 0 0100
   35 0010 + 0011 = 0 0101
   36 0010 + 0100 = 0 0110
   37 0010 + 0101 = 0 0111
   38 0010 + 0110 = 0 1000
   39 0010 + 0111 = 0 1001
   40 0010 + 1000 = 0 1010
   41 0010 + 1001 = 0 1011
   42 0010 + 1010 = 0 1100
   43 0010 + 1011 = 0 1101
   44 0010 + 1100 = 0 1110
   45 0010 + 1101 = 0 1111
   46 0010 + 1110 = 1 0000
   47 0010 + 1111 = 1 0001
   48 0011 + 0000 = 0 0011
   49 0011 + 0001 = 0 0100
   50 0011 + 0010 = 0 0101
   51 0011 + 0011 = 0 0110
   52 0011 + 0100 = 0 0111
   53 0011 + 0101 = 0 1000
   54 0011 + 0110 = 0 1001
   55 0011 + 0111 = 0 1010
   56 0011 + 1000 = 0 1011
   57 0011 + 1001 = 0 1100
   58 0011 + 1010 = 0 1101
   59 0011 + 1011 = 0 1110
   60 0011 + 1100 = 0 1111
   61 0011 + 1101 = 1 0000
   62 0011 + 1110 = 1 0001
   63 0011 + 1111 = 1 0010
   64 0100 + 0000 = 0 0100
   65 0100 + 0001 = 0 0101
   66 0100 + 0010 = 0 0110
   67 0100 + 0011 = 0 0111
   68 0100 + 0100 = 0 1000
   69 0100 + 0101 = 0 1001
   70 0100 + 0110 = 0 1010
   71 0100 + 0111 = 0 1011
   72 0100 + 1000 = 0 1100
   73 0100 + 1001 = 0 1101
   74 0100 + 1010 = 0 1110
   75 0100 + 1011 = 0 1111
   76 0100 + 1100 = 1 0000
   77 0100 + 1101 = 1 0001
   78 0100 + 1110 = 1 0010
   79 0100 + 1111 = 1 0011
   80 0101 + 0000 = 0 0101
   81 0101 + 0001 = 0 0110
   82 0101 + 0010 = 0 0111
   83 0101 + 0011 = 0 1000
   84 0101 + 0100 = 0 1001
   85 0101 + 0101 = 0 1010
   86 0101 + 0110 = 0 1011
   87 0101 + 0111 = 0 1100
   88 0101 + 1000 = 0 1101
   89 0101 + 1001 = 0 1110
   90 0101 + 1010 = 0 1111
   91 0101 + 1011 = 1 0000
   92 0101 + 1100 = 1 0001
   93 0101 + 1101 = 1 0010
   94 0101 + 1110 = 1 0011
   95 0101 + 1111 = 1 0100
   96 0110 + 0000 = 0 0110
   97 0110 + 0001 = 0 0111
   98 0110 + 0010 = 0 1000
   99 0110 + 0011 = 0 1001
  100 0110 + 0100 = 0 1010
  101 0110 + 0101 = 0 1011
  102 0110 + 0110 = 0 1100
  103 0110 + 0111 = 0 1101
  104 0110 + 1000 = 0 1110
  105 0110 + 1001 = 0 1111
  106 0110 + 1010 = 1 0000
  107 0110 + 1011 = 1 0001
  108 0110 + 1100 = 1 0010
  109 0110 + 1101 = 1 0011
  110 0110 + 1110 = 1 0100
  111 0110 + 1111 = 1 0101
  112 0111 + 0000 = 0 0111
  113 0111 + 0001 = 0 1000
  114 0111 + 0010 = 0 1001
  115 0111 + 0011 = 0 1010
  116 0111 + 0100 = 0 1011
  117 0111 + 0101 = 0 1100
  118 0111 + 0110 = 0 1101
  119 0111 + 0111 = 0 1110
  120 0111 + 1000 = 0 1111
  121 0111 + 1001 = 1 0000
  122 0111 + 1010 = 1 0001
  123 0111 + 1011 = 1 0010
  124 0111 + 1100 = 1 0011
  125 0111 + 1101 = 1 0100
  126 0111 + 1110 = 1 0101
  127 0111 + 1111 = 1 0110
  128 1000 + 0000 = 0 1000
  129 1000 + 0001 = 0 1001
  130 1000 + 0010 = 0 1010
  131 1000 + 0011 = 0 1011
  132 1000 + 0100 = 0 1100
  133 1000 + 0101 = 0 1101
  134 1000 + 0110 = 0 1110
  135 1000 + 0111 = 0 1111
  136 1000 + 1000 = 1 0000
  137 1000 + 1001 = 1 0001
  138 1000 + 1010 = 1 0010
  139 1000 + 1011 = 1 0011
  140 1000 + 1100 = 1 0100
  141 1000 + 1101 = 1 0101
  142 1000 + 1110 = 1 0110
  143 1000 + 1111 = 1 0111
  144 1001 + 0000 = 0 1001
  145 1001 + 0001 = 0 1010
  146 1001 + 0010 = 0 1011
  147 1001 + 0011 = 0 1100
  148 1001 + 0100 = 0 1101
  149 1001 + 0101 = 0 1110
  150 1001 + 0110 = 0 1111
  151 1001 + 0111 = 1 0000
  152 1001 + 1000 = 1 0001
  153 1001 + 1001 = 1 0010
  154 1001 + 1010 = 1 0011
  155 1001 + 1011 = 1 0100
  156 1001 + 1100 = 1 0101
  157 1001 + 1101 = 1 0110
  158 1001 + 1110 = 1 0111
  159 1001 + 1111 = 1 1000
  160 1010 + 0000 = 0 1010
  161 1010 + 0001 = 0 1011
  162 1010 + 0010 = 0 1100
  163 1010 + 0011 = 0 1101
  164 1010 + 0100 = 0 1110
  165 1010 + 0101 = 0 1111
  166 1010 + 0110 = 1 0000
  167 1010 + 0111 = 1 0001
  168 1010 + 1000 = 1 0010
  169 1010 + 1001 = 1 0011
  170 1010 + 1010 = 1 0100
  171 1010 + 1011 = 1 0101
  172 1010 + 1100 = 1 0110
  173 1010 + 1101 = 1 0111
  174 1010 + 1110 = 1 1000
  175 1010 + 1111 = 1 1001
  176 1011 + 0000 = 0 1011
  177 1011 + 0001 = 0 1100
  178 1011 + 0010 = 0 1101
  179 1011 + 0011 = 0 1110
  180 1011 + 0100 = 0 1111
  181 1011 + 0101 = 1 0000
  182 1011 + 0110 = 1 0001
  183 1011 + 0111 = 1 0010
  184 1011 + 1000 = 1 0011
  185 1011 + 1001 = 1 0100
  186 1011 + 1010 = 1 0101
  187 1011 + 1011 = 1 0110
  188 1011 + 1100 = 1 0111
  189 1011 + 1101 = 1 1000
  190 1011 + 1110 = 1 1001
  191 1011 + 1111 = 1 1010
  192 1100 + 0000 = 0 1100
  193 1100 + 0001 = 0 1101
  194 1100 + 0010 = 0 1110
  195 1100 + 0011 = 0 1111
  196 1100 + 0100 = 1 0000
  197 1100 + 0101 = 1 0001
  198 1100 + 0110 = 1 0010
  199 1100 + 0111 = 1 0011
  200 1100 + 1000 = 1 0100
  201 1100 + 1001 = 1 0101
  202 1100 + 1010 = 1 0110
  203 1100 + 1011 = 1 0111
  204 1100 + 1100 = 1 1000
  205 1100 + 1101 = 1 1001
  206 1100 + 1110 = 1 1010
  207 1100 + 1111 = 1 1011
  208 1101 + 0000 = 0 1101
  209 1101 + 0001 = 0 1110
  210 1101 + 0010 = 0 1111
  211 1101 + 0011 = 1 0000
  212 1101 + 0100 = 1 0001
  213 1101 + 0101 = 1 0010
  214 1101 + 0110 = 1 0011
  215 1101 + 0111 = 1 0100
  216 1101 + 1000 = 1 0101
  217 1101 + 1001 = 1 0110
  218 1101 + 1010 = 1 0111
  219 1101 + 1011 = 1 1000
  220 1101 + 1100 = 1 1001
  221 1101 + 1101 = 1 1010
  222 1101 + 1110 = 1 1011
  223 1101 + 1111 = 1 1100
  224 1110 + 0000 = 0 1110
  225 1110 + 0001 = 0 1111
  226 1110 + 0010 = 1 0000
  227 1110 + 0011 = 1 0001
  228 1110 + 0100 = 1 0010
  229 1110 + 0101 = 1 0011
  230 1110 + 0110 = 1 0100
  231 1110 + 0111 = 1 0101
  232 1110 + 1000 = 1 0110
  233 1110 + 1001 = 1 0111
  234 1110 + 1010 = 1 1000
  235 1110 + 1011 = 1 1001
  236 1110 + 1100 = 1 1010
  237 1110 + 1101 = 1 1011
  238 1110 + 1110 = 1 1100
  239 1110 + 1111 = 1 1101
  240 1111 + 0000 = 0 1111
  241 1111 + 0001 = 1 0000
  242 1111 + 0010 = 1 0001
  243 1111 + 0011 = 1 0010
  244 1111 + 0100 = 1 0011
  245 1111 + 0101 = 1 0100
  246 1111 + 0110 = 1 0101
  247 1111 + 0111 = 1 0110
  248 1111 + 1000 = 1 0111
  249 1111 + 1001 = 1 1000
  250 1111 + 1010 = 1 1001
  251 1111 + 1011 = 1 1010
  252 1111 + 1100 = 1 1011
  253 1111 + 1101 = 1 1100
  254 1111 + 1110 = 1 1101
  255 1111 + 1111 = 1 1110
*/

endmodule

