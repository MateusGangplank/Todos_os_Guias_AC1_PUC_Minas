// -----------------------------------------------------
// Guia 06_03 - Somador subtrator 4 bits compl 1
// Nome: Ludmily Caldeira da Silva
// Matricula: 417290
// -----------------------------------------------------

// -------------------------------------------------
// -- Somador subtrator 4 bits compl 1
// -------------------------------------------------

module MS (Soma, Cout, x, y);

output Cout, Soma;
input x, y;

xor XOR1 (Soma, x, y);
and AND1 (Cout, x, y);

endmodule // MS

module SC (Soma1, Cout1, x1, y1, Cin);

output Cout1, Soma1;
input x1, y1, Cin;
wire t1, t2, t3;

MS MS1 (t2, t1, x1, y1);
MS MS2 (Soma1, t3, Cin, t2);
or Or1 (Cout1, t3, t1);

endmodule // SC

module compLogico (s, a, b);

output s;
input [3:0]a;
input [3:0]b;
wire t1, t2, t3, t4;

xnor XNOR1 (t1, a[0], b[0]);
xnor XNOR2 (t2, a[1], b[1]);
xnor XNOR3 (t3, a[2], b[2]);
xnor XNOR4 (t4, a[3], b[3]);
and AND1 (s, t1, t2, t3, t4);

endmodule // compLogico

module compAritmetico (menor, maior, a, b);

output menor, maior;
input [3:0]a;
input [3:0]b;
wire t[0:7];
wire t1, t2, t3, t4;


xnor XNOR2 (t2, a[1], b[1]);
xnor XNOR3 (t3, a[2], b[2]);
xnor XNOR4 (t4, a[3], b[3]);

and AND1 (t[0], a[0], ~b[0], t4, t3, t2);
and AND2 (t[1], a[1], ~b[1], t4, t3);
and AND3 (t[2], a[2], ~b[2], t4);
and AND4 (t[3], a[3], ~b[3]);

or OR1 (maior, t[0], t[1], t[2], t[3]);

and AND5 (t[4], ~a[0], b[0], t4, t3, t2);
and AND6 (t[5], ~a[1], b[1], t4, t3);
and AND7 (t[6], ~a[2], b[2], t4);
and AND8 (t[7], ~a[3], b[3]);

or OR2 (menor, t[4], t[5], t[6], t[7]);

endmodule // compAritmetico


module SomaSubLogAriDetCompl (compl ,s2 ,maior, menor, s1, s, vout, a, b, sel);

output vout, s1, maior, menor, s2; 
output [3:0]s;
output [3:0]compl;
input sel;
input [3:0]a;
input [3:0]b; 
wire v[0:6];

xor XOR1 (v[0], sel, b[0]);
xor XOR2 (v[1], sel, b[1]);
xor XOR3 (v[2], sel, b[2]);
xor XOR4 (v[3], sel, b[3]);

SC SC0 (s[0], v[4], a[0], v[0], sel);
SC SC1 (s[1], v[5], a[1], v[1], v[4]);
SC SC2 (s[2], v[6], a[2], v[2], v[5]);
SC SC3 (s[3], vout, a[3], v[3], v[6]);

and AND1 (s2, sel, ~vout);

not Not2 (compl[0], s[0]);
not Not3 (compl[1], s[1]);
not Not4 (compl[2], s[2]);
not Not5 (compl[3], s[3]);

compLogico compLogico1 (s1, a, b);

compAritmetico CA (menor, maior, a, b);

endmodule // SomaSubLogAriDet

// -------------------------------------------------
// -- test Somador subtrator 4 bits compl 1
// -------------------------------------------------

module testSomaSubLogAriDetCompl;

reg [3:0]x;
reg [3:0]y;
reg sel;
wire [3:0]s;
wire [3:0]s3;
wire s1, s2;
wire cout, maior, menor;
integer j, k;

// instancia 
SomaSubLogAriDetCompl COMPL1 (s3, s2 ,maior, menor, s1, s, cout, x, y, sel);

// parte principal

initial begin
sel = 0;
x = 0;
y = 0;
j = 0;

end

 initial begin 
 
      $display("\nguia06_04 - Ludmily Caldeira da Silva - 417290\n");
      $display("Test Somador Completo 4 bits com comparador logico e aritmetico, detector e complemento de 1\n");      
		$display("\nSel    a      b      Cout  Soma/Subt   Compl 1   a = b      a > b   a < b  detector\n");
      $monitor("%b     %4b    %4b     %b     %4b       %4b       %b          %b       %b       %b" , sel, x, y, cout, s, s3, s1, maior, menor, s2);
		
		for (j = 0; j < 16; j = j + 1) begin
					
			#1 x = j;		
													
				for (k = 0; k < 16; k = k + 1) begin
		
					#1 y = k; 					
								
			   end
				
		   end
					
			for (j = 0; j < 16; j = j + 1) begin
					
			#1 x = j; sel = 1;
													
				for (k = 0; k < 16; k = k + 1) begin
		
					#1 y = k; 					
								
			   end
		
	   end		
				
  end
 
endmodule // testSomaSubLogAridetCompl 

/* Resultados obtidos
     
    
     ----jGRASP exec: vvp guia06-04.vvp
    
    
    guia06_04 - Ludmily Caldeira da Silva - 417290
    
    Test Somador Completo 4 bits com comparador logico e aritmetico, detector e complemento de 1
    
    
    Sel    a      b      Cout  Soma/Subt   Compl 1   a = b      a > b   a < b  detector
    
    0     0000    0000     0     0000       1111       1          0       0       0
    0     0000    0001     0     0001       1110       0          0       1       0
    0     0000    0010     0     0010       1101       0          0       1       0
    0     0000    0011     0     0011       1100       0          0       1       0
    0     0000    0100     0     0100       1011       0          0       1       0
    0     0000    0101     0     0101       1010       0          0       1       0
    0     0000    0110     0     0110       1001       0          0       1       0
    0     0000    0111     0     0111       1000       0          0       1       0
    0     0000    1000     0     1000       0111       0          0       1       0
    0     0000    1001     0     1001       0110       0          0       1       0
    0     0000    1010     0     1010       0101       0          0       1       0
    0     0000    1011     0     1011       0100       0          0       1       0
    0     0000    1100     0     1100       0011       0          0       1       0
    0     0000    1101     0     1101       0010       0          0       1       0
    0     0000    1110     0     1110       0001       0          0       1       0
    0     0000    1111     0     1111       0000       0          0       1       0
    0     0001    1111     1     0000       1111       0          0       1       0
    0     0001    0000     0     0001       1110       0          1       0       0
    0     0001    0001     0     0010       1101       1          0       0       0
    0     0001    0010     0     0011       1100       0          0       1       0
    0     0001    0011     0     0100       1011       0          0       1       0
    0     0001    0100     0     0101       1010       0          0       1       0
    0     0001    0101     0     0110       1001       0          0       1       0
    0     0001    0110     0     0111       1000       0          0       1       0
    0     0001    0111     0     1000       0111       0          0       1       0
    0     0001    1000     0     1001       0110       0          0       1       0
    0     0001    1001     0     1010       0101       0          0       1       0
    0     0001    1010     0     1011       0100       0          0       1       0
    0     0001    1011     0     1100       0011       0          0       1       0
    0     0001    1100     0     1101       0010       0          0       1       0
    0     0001    1101     0     1110       0001       0          0       1       0
    0     0001    1110     0     1111       0000       0          0       1       0
    0     0001    1111     1     0000       1111       0          0       1       0
    0     0010    1111     1     0001       1110       0          0       1       0
    0     0010    0000     0     0010       1101       0          1       0       0
    0     0010    0001     0     0011       1100       0          1       0       0
    0     0010    0010     0     0100       1011       1          0       0       0
    0     0010    0011     0     0101       1010       0          0       1       0
    0     0010    0100     0     0110       1001       0          0       1       0
    0     0010    0101     0     0111       1000       0          0       1       0
    0     0010    0110     0     1000       0111       0          0       1       0
    0     0010    0111     0     1001       0110       0          0       1       0
    0     0010    1000     0     1010       0101       0          0       1       0
    0     0010    1001     0     1011       0100       0          0       1       0
    0     0010    1010     0     1100       0011       0          0       1       0
    0     0010    1011     0     1101       0010       0          0       1       0
    0     0010    1100     0     1110       0001       0          0       1       0
    0     0010    1101     0     1111       0000       0          0       1       0
    0     0010    1110     1     0000       1111       0          0       1       0
    0     0010    1111     1     0001       1110       0          0       1       0
    0     0011    1111     1     0010       1101       0          0       1       0
    0     0011    0000     0     0011       1100       0          1       0       0
    0     0011    0001     0     0100       1011       0          1       0       0
    0     0011    0010     0     0101       1010       0          1       0       0
    0     0011    0011     0     0110       1001       1          0       0       0
    0     0011    0100     0     0111       1000       0          0       1       0
    0     0011    0101     0     1000       0111       0          0       1       0
    0     0011    0110     0     1001       0110       0          0       1       0
    0     0011    0111     0     1010       0101       0          0       1       0
    0     0011    1000     0     1011       0100       0          0       1       0
    0     0011    1001     0     1100       0011       0          0       1       0
    0     0011    1010     0     1101       0010       0          0       1       0
    0     0011    1011     0     1110       0001       0          0       1       0
    0     0011    1100     0     1111       0000       0          0       1       0
    0     0011    1101     1     0000       1111       0          0       1       0
    0     0011    1110     1     0001       1110       0          0       1       0
    0     0011    1111     1     0010       1101       0          0       1       0
    0     0100    1111     1     0011       1100       0          0       1       0
    0     0100    0000     0     0100       1011       0          1       0       0
    0     0100    0001     0     0101       1010       0          1       0       0
    0     0100    0010     0     0110       1001       0          1       0       0
    0     0100    0011     0     0111       1000       0          1       0       0
    0     0100    0100     0     1000       0111       1          0       0       0
    0     0100    0101     0     1001       0110       0          0       1       0
    0     0100    0110     0     1010       0101       0          0       1       0
    0     0100    0111     0     1011       0100       0          0       1       0
    0     0100    1000     0     1100       0011       0          0       1       0
    0     0100    1001     0     1101       0010       0          0       1       0
    0     0100    1010     0     1110       0001       0          0       1       0
    0     0100    1011     0     1111       0000       0          0       1       0
    0     0100    1100     1     0000       1111       0          0       1       0
    0     0100    1101     1     0001       1110       0          0       1       0
    0     0100    1110     1     0010       1101       0          0       1       0
    0     0100    1111     1     0011       1100       0          0       1       0
    0     0101    1111     1     0100       1011       0          0       1       0
    0     0101    0000     0     0101       1010       0          1       0       0
    0     0101    0001     0     0110       1001       0          1       0       0
    0     0101    0010     0     0111       1000       0          1       0       0
    0     0101    0011     0     1000       0111       0          1       0       0
    0     0101    0100     0     1001       0110       0          1       0       0
    0     0101    0101     0     1010       0101       1          0       0       0
    0     0101    0110     0     1011       0100       0          0       1       0
    0     0101    0111     0     1100       0011       0          0       1       0
    0     0101    1000     0     1101       0010       0          0       1       0
    0     0101    1001     0     1110       0001       0          0       1       0
    0     0101    1010     0     1111       0000       0          0       1       0
    0     0101    1011     1     0000       1111       0          0       1       0
    0     0101    1100     1     0001       1110       0          0       1       0
    0     0101    1101     1     0010       1101       0          0       1       0
    0     0101    1110     1     0011       1100       0          0       1       0
    0     0101    1111     1     0100       1011       0          0       1       0
    0     0110    1111     1     0101       1010       0          0       1       0
    0     0110    0000     0     0110       1001       0          1       0       0
    0     0110    0001     0     0111       1000       0          1       0       0
    0     0110    0010     0     1000       0111       0          1       0       0
    0     0110    0011     0     1001       0110       0          1       0       0
    0     0110    0100     0     1010       0101       0          1       0       0
    0     0110    0101     0     1011       0100       0          1       0       0
    0     0110    0110     0     1100       0011       1          0       0       0
    0     0110    0111     0     1101       0010       0          0       1       0
    0     0110    1000     0     1110       0001       0          0       1       0
    0     0110    1001     0     1111       0000       0          0       1       0
    0     0110    1010     1     0000       1111       0          0       1       0
    0     0110    1011     1     0001       1110       0          0       1       0
    0     0110    1100     1     0010       1101       0          0       1       0
    0     0110    1101     1     0011       1100       0          0       1       0
    0     0110    1110     1     0100       1011       0          0       1       0
    0     0110    1111     1     0101       1010       0          0       1       0
    0     0111    1111     1     0110       1001       0          0       1       0
    0     0111    0000     0     0111       1000       0          1       0       0
    0     0111    0001     0     1000       0111       0          1       0       0
    0     0111    0010     0     1001       0110       0          1       0       0
    0     0111    0011     0     1010       0101       0          1       0       0
    0     0111    0100     0     1011       0100       0          1       0       0
    0     0111    0101     0     1100       0011       0          1       0       0
    0     0111    0110     0     1101       0010       0          1       0       0
    0     0111    0111     0     1110       0001       1          0       0       0
    0     0111    1000     0     1111       0000       0          0       1       0
    0     0111    1001     1     0000       1111       0          0       1       0
    0     0111    1010     1     0001       1110       0          0       1       0
    0     0111    1011     1     0010       1101       0          0       1       0
    0     0111    1100     1     0011       1100       0          0       1       0
    0     0111    1101     1     0100       1011       0          0       1       0
    0     0111    1110     1     0101       1010       0          0       1       0
    0     0111    1111     1     0110       1001       0          0       1       0
    0     1000    1111     1     0111       1000       0          0       1       0
    0     1000    0000     0     1000       0111       0          1       0       0
    0     1000    0001     0     1001       0110       0          1       0       0
    0     1000    0010     0     1010       0101       0          1       0       0
    0     1000    0011     0     1011       0100       0          1       0       0
    0     1000    0100     0     1100       0011       0          1       0       0
    0     1000    0101     0     1101       0010       0          1       0       0
    0     1000    0110     0     1110       0001       0          1       0       0
    0     1000    0111     0     1111       0000       0          1       0       0
    0     1000    1000     1     0000       1111       1          0       0       0
    0     1000    1001     1     0001       1110       0          0       1       0
    0     1000    1010     1     0010       1101       0          0       1       0
    0     1000    1011     1     0011       1100       0          0       1       0
    0     1000    1100     1     0100       1011       0          0       1       0
    0     1000    1101     1     0101       1010       0          0       1       0
    0     1000    1110     1     0110       1001       0          0       1       0
    0     1000    1111     1     0111       1000       0          0       1       0
    0     1001    1111     1     1000       0111       0          0       1       0
    0     1001    0000     0     1001       0110       0          1       0       0
    0     1001    0001     0     1010       0101       0          1       0       0
    0     1001    0010     0     1011       0100       0          1       0       0
    0     1001    0011     0     1100       0011       0          1       0       0
    0     1001    0100     0     1101       0010       0          1       0       0
    0     1001    0101     0     1110       0001       0          1       0       0
    0     1001    0110     0     1111       0000       0          1       0       0
    0     1001    0111     1     0000       1111       0          1       0       0
    0     1001    1000     1     0001       1110       0          1       0       0
    0     1001    1001     1     0010       1101       1          0       0       0
    0     1001    1010     1     0011       1100       0          0       1       0
    0     1001    1011     1     0100       1011       0          0       1       0
    0     1001    1100     1     0101       1010       0          0       1       0
    0     1001    1101     1     0110       1001       0          0       1       0
    0     1001    1110     1     0111       1000       0          0       1       0
    0     1001    1111     1     1000       0111       0          0       1       0
    0     1010    1111     1     1001       0110       0          0       1       0
    0     1010    0000     0     1010       0101       0          1       0       0
    0     1010    0001     0     1011       0100       0          1       0       0
    0     1010    0010     0     1100       0011       0          1       0       0
    0     1010    0011     0     1101       0010       0          1       0       0
    0     1010    0100     0     1110       0001       0          1       0       0
    0     1010    0101     0     1111       0000       0          1       0       0
    0     1010    0110     1     0000       1111       0          1       0       0
    0     1010    0111     1     0001       1110       0          1       0       0
    0     1010    1000     1     0010       1101       0          1       0       0
    0     1010    1001     1     0011       1100       0          1       0       0
    0     1010    1010     1     0100       1011       1          0       0       0
    0     1010    1011     1     0101       1010       0          0       1       0
    0     1010    1100     1     0110       1001       0          0       1       0
    0     1010    1101     1     0111       1000       0          0       1       0
    0     1010    1110     1     1000       0111       0          0       1       0
    0     1010    1111     1     1001       0110       0          0       1       0
    0     1011    1111     1     1010       0101       0          0       1       0
    0     1011    0000     0     1011       0100       0          1       0       0
    0     1011    0001     0     1100       0011       0          1       0       0
    0     1011    0010     0     1101       0010       0          1       0       0
    0     1011    0011     0     1110       0001       0          1       0       0
    0     1011    0100     0     1111       0000       0          1       0       0
    0     1011    0101     1     0000       1111       0          1       0       0
    0     1011    0110     1     0001       1110       0          1       0       0
    0     1011    0111     1     0010       1101       0          1       0       0
    0     1011    1000     1     0011       1100       0          1       0       0
    0     1011    1001     1     0100       1011       0          1       0       0
    0     1011    1010     1     0101       1010       0          1       0       0
    0     1011    1011     1     0110       1001       1          0       0       0
    0     1011    1100     1     0111       1000       0          0       1       0
    0     1011    1101     1     1000       0111       0          0       1       0
    0     1011    1110     1     1001       0110       0          0       1       0
    0     1011    1111     1     1010       0101       0          0       1       0
    0     1100    1111     1     1011       0100       0          0       1       0
    0     1100    0000     0     1100       0011       0          1       0       0
    0     1100    0001     0     1101       0010       0          1       0       0
    0     1100    0010     0     1110       0001       0          1       0       0
    0     1100    0011     0     1111       0000       0          1       0       0
    0     1100    0100     1     0000       1111       0          1       0       0
    0     1100    0101     1     0001       1110       0          1       0       0
    0     1100    0110     1     0010       1101       0          1       0       0
    0     1100    0111     1     0011       1100       0          1       0       0
    0     1100    1000     1     0100       1011       0          1       0       0
    0     1100    1001     1     0101       1010       0          1       0       0
    0     1100    1010     1     0110       1001       0          1       0       0
    0     1100    1011     1     0111       1000       0          1       0       0
    0     1100    1100     1     1000       0111       1          0       0       0
    0     1100    1101     1     1001       0110       0          0       1       0
    0     1100    1110     1     1010       0101       0          0       1       0
    0     1100    1111     1     1011       0100       0          0       1       0
    0     1101    1111     1     1100       0011       0          0       1       0
    0     1101    0000     0     1101       0010       0          1       0       0
    0     1101    0001     0     1110       0001       0          1       0       0
    0     1101    0010     0     1111       0000       0          1       0       0
    0     1101    0011     1     0000       1111       0          1       0       0
    0     1101    0100     1     0001       1110       0          1       0       0
    0     1101    0101     1     0010       1101       0          1       0       0
    0     1101    0110     1     0011       1100       0          1       0       0
    0     1101    0111     1     0100       1011       0          1       0       0
    0     1101    1000     1     0101       1010       0          1       0       0
    0     1101    1001     1     0110       1001       0          1       0       0
    0     1101    1010     1     0111       1000       0          1       0       0
    0     1101    1011     1     1000       0111       0          1       0       0
    0     1101    1100     1     1001       0110       0          1       0       0
    0     1101    1101     1     1010       0101       1          0       0       0
    0     1101    1110     1     1011       0100       0          0       1       0
    0     1101    1111     1     1100       0011       0          0       1       0
    0     1110    1111     1     1101       0010       0          0       1       0
    0     1110    0000     0     1110       0001       0          1       0       0
    0     1110    0001     0     1111       0000       0          1       0       0
    0     1110    0010     1     0000       1111       0          1       0       0
    0     1110    0011     1     0001       1110       0          1       0       0
    0     1110    0100     1     0010       1101       0          1       0       0
    0     1110    0101     1     0011       1100       0          1       0       0
    0     1110    0110     1     0100       1011       0          1       0       0
    0     1110    0111     1     0101       1010       0          1       0       0
    0     1110    1000     1     0110       1001       0          1       0       0
    0     1110    1001     1     0111       1000       0          1       0       0
    0     1110    1010     1     1000       0111       0          1       0       0
    0     1110    1011     1     1001       0110       0          1       0       0
    0     1110    1100     1     1010       0101       0          1       0       0
    0     1110    1101     1     1011       0100       0          1       0       0
    0     1110    1110     1     1100       0011       1          0       0       0
    0     1110    1111     1     1101       0010       0          0       1       0
    0     1111    1111     1     1110       0001       1          0       0       0
    0     1111    0000     0     1111       0000       0          1       0       0
    0     1111    0001     1     0000       1111       0          1       0       0
    0     1111    0010     1     0001       1110       0          1       0       0
    0     1111    0011     1     0010       1101       0          1       0       0
    0     1111    0100     1     0011       1100       0          1       0       0
    0     1111    0101     1     0100       1011       0          1       0       0
    0     1111    0110     1     0101       1010       0          1       0       0
    0     1111    0111     1     0110       1001       0          1       0       0
    0     1111    1000     1     0111       1000       0          1       0       0
    0     1111    1001     1     1000       0111       0          1       0       0
    0     1111    1010     1     1001       0110       0          1       0       0
    0     1111    1011     1     1010       0101       0          1       0       0
    0     1111    1100     1     1011       0100       0          1       0       0
    0     1111    1101     1     1100       0011       0          1       0       0
    0     1111    1110     1     1101       0010       0          1       0       0
    0     1111    1111     1     1110       0001       1          0       0       0
    1     0000    1111     0     0001       1110       0          0       1       1
    1     0000    0000     1     0000       1111       1          0       0       0
    1     0000    0001     0     1111       0000       0          0       1       1
    1     0000    0010     0     1110       0001       0          0       1       1
    1     0000    0011     0     1101       0010       0          0       1       1
    1     0000    0100     0     1100       0011       0          0       1       1
    1     0000    0101     0     1011       0100       0          0       1       1
    1     0000    0110     0     1010       0101       0          0       1       1
    1     0000    0111     0     1001       0110       0          0       1       1
    1     0000    1000     0     1000       0111       0          0       1       1
    1     0000    1001     0     0111       1000       0          0       1       1
    1     0000    1010     0     0110       1001       0          0       1       1
    1     0000    1011     0     0101       1010       0          0       1       1
    1     0000    1100     0     0100       1011       0          0       1       1
    1     0000    1101     0     0011       1100       0          0       1       1
    1     0000    1110     0     0010       1101       0          0       1       1
    1     0000    1111     0     0001       1110       0          0       1       1
    1     0001    1111     0     0010       1101       0          0       1       1
    1     0001    0000     1     0001       1110       0          1       0       0
    1     0001    0001     1     0000       1111       1          0       0       0
    1     0001    0010     0     1111       0000       0          0       1       1
    1     0001    0011     0     1110       0001       0          0       1       1
    1     0001    0100     0     1101       0010       0          0       1       1
    1     0001    0101     0     1100       0011       0          0       1       1
    1     0001    0110     0     1011       0100       0          0       1       1
    1     0001    0111     0     1010       0101       0          0       1       1
    1     0001    1000     0     1001       0110       0          0       1       1
    1     0001    1001     0     1000       0111       0          0       1       1
    1     0001    1010     0     0111       1000       0          0       1       1
    1     0001    1011     0     0110       1001       0          0       1       1
    1     0001    1100     0     0101       1010       0          0       1       1
    1     0001    1101     0     0100       1011       0          0       1       1
    1     0001    1110     0     0011       1100       0          0       1       1
    1     0001    1111     0     0010       1101       0          0       1       1
    1     0010    1111     0     0011       1100       0          0       1       1
    1     0010    0000     1     0010       1101       0          1       0       0
    1     0010    0001     1     0001       1110       0          1       0       0
    1     0010    0010     1     0000       1111       1          0       0       0
    1     0010    0011     0     1111       0000       0          0       1       1
    1     0010    0100     0     1110       0001       0          0       1       1
    1     0010    0101     0     1101       0010       0          0       1       1
    1     0010    0110     0     1100       0011       0          0       1       1
    1     0010    0111     0     1011       0100       0          0       1       1
    1     0010    1000     0     1010       0101       0          0       1       1
    1     0010    1001     0     1001       0110       0          0       1       1
    1     0010    1010     0     1000       0111       0          0       1       1
    1     0010    1011     0     0111       1000       0          0       1       1
    1     0010    1100     0     0110       1001       0          0       1       1
    1     0010    1101     0     0101       1010       0          0       1       1
    1     0010    1110     0     0100       1011       0          0       1       1
    1     0010    1111     0     0011       1100       0          0       1       1
    1     0011    1111     0     0100       1011       0          0       1       1
    1     0011    0000     1     0011       1100       0          1       0       0
    1     0011    0001     1     0010       1101       0          1       0       0
    1     0011    0010     1     0001       1110       0          1       0       0
    1     0011    0011     1     0000       1111       1          0       0       0
    1     0011    0100     0     1111       0000       0          0       1       1
    1     0011    0101     0     1110       0001       0          0       1       1
    1     0011    0110     0     1101       0010       0          0       1       1
    1     0011    0111     0     1100       0011       0          0       1       1
    1     0011    1000     0     1011       0100       0          0       1       1
    1     0011    1001     0     1010       0101       0          0       1       1
    1     0011    1010     0     1001       0110       0          0       1       1
    1     0011    1011     0     1000       0111       0          0       1       1
    1     0011    1100     0     0111       1000       0          0       1       1
    1     0011    1101     0     0110       1001       0          0       1       1
    1     0011    1110     0     0101       1010       0          0       1       1
    1     0011    1111     0     0100       1011       0          0       1       1
    1     0100    1111     0     0101       1010       0          0       1       1
    1     0100    0000     1     0100       1011       0          1       0       0
    1     0100    0001     1     0011       1100       0          1       0       0
    1     0100    0010     1     0010       1101       0          1       0       0
    1     0100    0011     1     0001       1110       0          1       0       0
    1     0100    0100     1     0000       1111       1          0       0       0
    1     0100    0101     0     1111       0000       0          0       1       1
    1     0100    0110     0     1110       0001       0          0       1       1
    1     0100    0111     0     1101       0010       0          0       1       1
    1     0100    1000     0     1100       0011       0          0       1       1
    1     0100    1001     0     1011       0100       0          0       1       1
    1     0100    1010     0     1010       0101       0          0       1       1
    1     0100    1011     0     1001       0110       0          0       1       1
    1     0100    1100     0     1000       0111       0          0       1       1
    1     0100    1101     0     0111       1000       0          0       1       1
    1     0100    1110     0     0110       1001       0          0       1       1
    1     0100    1111     0     0101       1010       0          0       1       1
    1     0101    1111     0     0110       1001       0          0       1       1
    1     0101    0000     1     0101       1010       0          1       0       0
    1     0101    0001     1     0100       1011       0          1       0       0
    1     0101    0010     1     0011       1100       0          1       0       0
    1     0101    0011     1     0010       1101       0          1       0       0
    1     0101    0100     1     0001       1110       0          1       0       0
    1     0101    0101     1     0000       1111       1          0       0       0
    1     0101    0110     0     1111       0000       0          0       1       1
    1     0101    0111     0     1110       0001       0          0       1       1
    1     0101    1000     0     1101       0010       0          0       1       1
    1     0101    1001     0     1100       0011       0          0       1       1
    1     0101    1010     0     1011       0100       0          0       1       1
    1     0101    1011     0     1010       0101       0          0       1       1
    1     0101    1100     0     1001       0110       0          0       1       1
    1     0101    1101     0     1000       0111       0          0       1       1
    1     0101    1110     0     0111       1000       0          0       1       1
    1     0101    1111     0     0110       1001       0          0       1       1
    1     0110    1111     0     0111       1000       0          0       1       1
    1     0110    0000     1     0110       1001       0          1       0       0
    1     0110    0001     1     0101       1010       0          1       0       0
    1     0110    0010     1     0100       1011       0          1       0       0
    1     0110    0011     1     0011       1100       0          1       0       0
    1     0110    0100     1     0010       1101       0          1       0       0
    1     0110    0101     1     0001       1110       0          1       0       0
    1     0110    0110     1     0000       1111       1          0       0       0
    1     0110    0111     0     1111       0000       0          0       1       1
    1     0110    1000     0     1110       0001       0          0       1       1
    1     0110    1001     0     1101       0010       0          0       1       1
    1     0110    1010     0     1100       0011       0          0       1       1
    1     0110    1011     0     1011       0100       0          0       1       1
    1     0110    1100     0     1010       0101       0          0       1       1
    1     0110    1101     0     1001       0110       0          0       1       1
    1     0110    1110     0     1000       0111       0          0       1       1
    1     0110    1111     0     0111       1000       0          0       1       1
    1     0111    1111     0     1000       0111       0          0       1       1
    1     0111    0000     1     0111       1000       0          1       0       0
    1     0111    0001     1     0110       1001       0          1       0       0
    1     0111    0010     1     0101       1010       0          1       0       0
    1     0111    0011     1     0100       1011       0          1       0       0
    1     0111    0100     1     0011       1100       0          1       0       0
    1     0111    0101     1     0010       1101       0          1       0       0
    1     0111    0110     1     0001       1110       0          1       0       0
    1     0111    0111     1     0000       1111       1          0       0       0
    1     0111    1000     0     1111       0000       0          0       1       1
    1     0111    1001     0     1110       0001       0          0       1       1
    1     0111    1010     0     1101       0010       0          0       1       1
    1     0111    1011     0     1100       0011       0          0       1       1
    1     0111    1100     0     1011       0100       0          0       1       1
    1     0111    1101     0     1010       0101       0          0       1       1
    1     0111    1110     0     1001       0110       0          0       1       1
    1     0111    1111     0     1000       0111       0          0       1       1
    1     1000    1111     0     1001       0110       0          0       1       1
    1     1000    0000     1     1000       0111       0          1       0       0
    1     1000    0001     1     0111       1000       0          1       0       0
    1     1000    0010     1     0110       1001       0          1       0       0
    1     1000    0011     1     0101       1010       0          1       0       0
    1     1000    0100     1     0100       1011       0          1       0       0
    1     1000    0101     1     0011       1100       0          1       0       0
    1     1000    0110     1     0010       1101       0          1       0       0
    1     1000    0111     1     0001       1110       0          1       0       0
    1     1000    1000     1     0000       1111       1          0       0       0
    1     1000    1001     0     1111       0000       0          0       1       1
    1     1000    1010     0     1110       0001       0          0       1       1
    1     1000    1011     0     1101       0010       0          0       1       1
    1     1000    1100     0     1100       0011       0          0       1       1
    1     1000    1101     0     1011       0100       0          0       1       1
    1     1000    1110     0     1010       0101       0          0       1       1
    1     1000    1111     0     1001       0110       0          0       1       1
    1     1001    1111     0     1010       0101       0          0       1       1
    1     1001    0000     1     1001       0110       0          1       0       0
    1     1001    0001     1     1000       0111       0          1       0       0
    1     1001    0010     1     0111       1000       0          1       0       0
    1     1001    0011     1     0110       1001       0          1       0       0
    1     1001    0100     1     0101       1010       0          1       0       0
    1     1001    0101     1     0100       1011       0          1       0       0
    1     1001    0110     1     0011       1100       0          1       0       0
    1     1001    0111     1     0010       1101       0          1       0       0
    1     1001    1000     1     0001       1110       0          1       0       0
    1     1001    1001     1     0000       1111       1          0       0       0
    1     1001    1010     0     1111       0000       0          0       1       1
    1     1001    1011     0     1110       0001       0          0       1       1
    1     1001    1100     0     1101       0010       0          0       1       1
    1     1001    1101     0     1100       0011       0          0       1       1
    1     1001    1110     0     1011       0100       0          0       1       1
    1     1001    1111     0     1010       0101       0          0       1       1
    1     1010    1111     0     1011       0100       0          0       1       1
    1     1010    0000     1     1010       0101       0          1       0       0
    1     1010    0001     1     1001       0110       0          1       0       0
    1     1010    0010     1     1000       0111       0          1       0       0
    1     1010    0011     1     0111       1000       0          1       0       0
    1     1010    0100     1     0110       1001       0          1       0       0
    1     1010    0101     1     0101       1010       0          1       0       0
    1     1010    0110     1     0100       1011       0          1       0       0
    1     1010    0111     1     0011       1100       0          1       0       0
    1     1010    1000     1     0010       1101       0          1       0       0
    1     1010    1001     1     0001       1110       0          1       0       0
    1     1010    1010     1     0000       1111       1          0       0       0
    1     1010    1011     0     1111       0000       0          0       1       1
    1     1010    1100     0     1110       0001       0          0       1       1
    1     1010    1101     0     1101       0010       0          0       1       1
    1     1010    1110     0     1100       0011       0          0       1       1
    1     1010    1111     0     1011       0100       0          0       1       1
    1     1011    1111     0     1100       0011       0          0       1       1
    1     1011    0000     1     1011       0100       0          1       0       0
    1     1011    0001     1     1010       0101       0          1       0       0
    1     1011    0010     1     1001       0110       0          1       0       0
    1     1011    0011     1     1000       0111       0          1       0       0
    1     1011    0100     1     0111       1000       0          1       0       0
    1     1011    0101     1     0110       1001       0          1       0       0
    1     1011    0110     1     0101       1010       0          1       0       0
    1     1011    0111     1     0100       1011       0          1       0       0
    1     1011    1000     1     0011       1100       0          1       0       0
    1     1011    1001     1     0010       1101       0          1       0       0
    1     1011    1010     1     0001       1110       0          1       0       0
    1     1011    1011     1     0000       1111       1          0       0       0
    1     1011    1100     0     1111       0000       0          0       1       1
    1     1011    1101     0     1110       0001       0          0       1       1
    1     1011    1110     0     1101       0010       0          0       1       1
    1     1011    1111     0     1100       0011       0          0       1       1
    1     1100    1111     0     1101       0010       0          0       1       1
    1     1100    0000     1     1100       0011       0          1       0       0
    1     1100    0001     1     1011       0100       0          1       0       0
    1     1100    0010     1     1010       0101       0          1       0       0
    1     1100    0011     1     1001       0110       0          1       0       0
    1     1100    0100     1     1000       0111       0          1       0       0
    1     1100    0101     1     0111       1000       0          1       0       0
    1     1100    0110     1     0110       1001       0          1       0       0
    1     1100    0111     1     0101       1010       0          1       0       0
    1     1100    1000     1     0100       1011       0          1       0       0
    1     1100    1001     1     0011       1100       0          1       0       0
    1     1100    1010     1     0010       1101       0          1       0       0
    1     1100    1011     1     0001       1110       0          1       0       0
    1     1100    1100     1     0000       1111       1          0       0       0
    1     1100    1101     0     1111       0000       0          0       1       1
    1     1100    1110     0     1110       0001       0          0       1       1
    1     1100    1111     0     1101       0010       0          0       1       1
    1     1101    1111     0     1110       0001       0          0       1       1
    1     1101    0000     1     1101       0010       0          1       0       0
    1     1101    0001     1     1100       0011       0          1       0       0
    1     1101    0010     1     1011       0100       0          1       0       0
    1     1101    0011     1     1010       0101       0          1       0       0
    1     1101    0100     1     1001       0110       0          1       0       0
    1     1101    0101     1     1000       0111       0          1       0       0
    1     1101    0110     1     0111       1000       0          1       0       0
    1     1101    0111     1     0110       1001       0          1       0       0
    1     1101    1000     1     0101       1010       0          1       0       0
    1     1101    1001     1     0100       1011       0          1       0       0
    1     1101    1010     1     0011       1100       0          1       0       0
    1     1101    1011     1     0010       1101       0          1       0       0
    1     1101    1100     1     0001       1110       0          1       0       0
    1     1101    1101     1     0000       1111       1          0       0       0
    1     1101    1110     0     1111       0000       0          0       1       1
    1     1101    1111     0     1110       0001       0          0       1       1
    1     1110    1111     0     1111       0000       0          0       1       1
    1     1110    0000     1     1110       0001       0          1       0       0
    1     1110    0001     1     1101       0010       0          1       0       0
    1     1110    0010     1     1100       0011       0          1       0       0
    1     1110    0011     1     1011       0100       0          1       0       0
    1     1110    0100     1     1010       0101       0          1       0       0
    1     1110    0101     1     1001       0110       0          1       0       0
    1     1110    0110     1     1000       0111       0          1       0       0
    1     1110    0111     1     0111       1000       0          1       0       0
    1     1110    1000     1     0110       1001       0          1       0       0
    1     1110    1001     1     0101       1010       0          1       0       0
    1     1110    1010     1     0100       1011       0          1       0       0
    1     1110    1011     1     0011       1100       0          1       0       0
    1     1110    1100     1     0010       1101       0          1       0       0
    1     1110    1101     1     0001       1110       0          1       0       0
    1     1110    1110     1     0000       1111       1          0       0       0
    1     1110    1111     0     1111       0000       0          0       1       1
    1     1111    1111     1     0000       1111       1          0       0       0
    1     1111    0000     1     1111       0000       0          1       0       0
    1     1111    0001     1     1110       0001       0          1       0       0
    1     1111    0010     1     1101       0010       0          1       0       0
    1     1111    0011     1     1100       0011       0          1       0       0
    1     1111    0100     1     1011       0100       0          1       0       0
    1     1111    0101     1     1010       0101       0          1       0       0
    1     1111    0110     1     1001       0110       0          1       0       0
    1     1111    0111     1     1000       0111       0          1       0       0
    1     1111    1000     1     0111       1000       0          1       0       0
    1     1111    1001     1     0110       1001       0          1       0       0
    1     1111    1010     1     0101       1010       0          1       0       0
    1     1111    1011     1     0100       1011       0          1       0       0
    1     1111    1100     1     0011       1100       0          1       0       0
    1     1111    1101     1     0010       1101       0          1       0       0
    1     1111    1110     1     0001       1110       0          1       0       0
    1     1111    1111     1     0000       1111       1          0       0       0
    
     ----jGRASP: operation complete.
             */