// ------------------------- 
// Exemplo0014 
// Nome: Miller 
// Matricula: 449048 
// ------------------------- 
 
// ------------------------- 
//  test number system 
// ------------------------- 
 
module test_base_04; 
// ------------------------- definir dados 
      reg [2:0] a; 
      reg [3:0] b; 
      reg [4:0] c; 
      reg [4:0] d; 
 
// ------------------------- parte principal 
 initial begin 
      $display("Exemplo0014 - Miller - 449048"); 
      $display("Test number system"); 
		
		a =   5; 
      b =  10; 
      c =  15; 
      d =  20; 
       
      $display("\nPositive value"); 
      $display("a = %d = %3b", a, a); 
      $display("b = %d = %4b", a, a); 
      $display("c = %d = %5b", a, a); 
 
      $display("b = %d = %4b", b, b); 
      $display("c = %d = %5b", c, c); 
      $display("d = %d = %5b", d, d); 
      $display("d = %d = %5o", d, d); 
      $display("d = %d = %5h", d, d);
		
		a = -5;
		b = -5;
		c = -5;
		$display("\nNegative value");
		$display("a = -5 [3] = %d = %3b", a, a);
		$display("b = -5 [4] = %d = %4b", b, b);
		$display("c = -5 [5] = %d = %5b", c, c);
 
      a = ~5+1; 
      b = ~5+1; 
      c = ~5+1; 
 
      $display("\nNegative mixed expression"); 
      $display("a = %d = %3b", a, a); 
      $display("b = %d = %4b", b, b); 
      $display("c = %d = %5b", c, c);
		
		a = 5 + 3; 
		b = 5 + 3; 
 		c = 10 - 5 + 25 + 3 + 1; 
 		$display("\nOverflow"); 
 		$display("a = %d = %3b", a, a); 
 		$display("b = %d = %4b", b, b); 
 		$display("c = %d = %5b", c, c); 
		
		end 
 
endmodule // test_base

//-- Obs.:
//-- Ficar de olho na quantidade de bits e aumentar em 1 ou 2 casas em caso de soma,
//-- para evitar um overflow, "espa�o insuficiente" !
//-- O tamanho de cada variavel ja foi definida no reg[x:0] la em cima, reprensentando o seu tamanho.
//-- reg [2:0] = 3 bits de representacao;
//-- reg [7:0] = 8 bits de representacao;
//-- por isso, quando colocamos %d utilizando a varivel a da 0, pois a variavel a, inicialmente possui
//-- 3 bits de representa�ao, reg [2:0] a; , e o 8 = 1000 , 4 bits, ou seja, apenas 000 foi armazenado.




