// ---------------------
// Guia 05_01 - 4 bits Full Adder with NOR gate
// Nome: Alyson Deives
// Matricula: 416589
// ---------------------

// -------------------------------
// -- 4 bits full adder with with NOR gate
// -------------------------------

module four_bits_fulladder_nor (c,a,b);
output [4:0] c;
input [3:0] a;
input [3:0] b;


halfadder_nor HA1 (c[0],carry1,a[0],b[0]);
fulladder_nor FA1 (c[1],carry2,a[1],b[1],carry1);
fulladder_nor FA2 (c[2],carry3,a[2],b[2],carry2);
fulladder_nor FA3 (c[3],c[4],a[3],b[3],carry3);

endmodule // 4_bits_full_adder_nor


// -------------------------------
// -- full adder with NOR gate
// -------------------------------

module fulladder_nor (c0,c1,r,s,t);
output c0,c1;
input r,s,t;
wire carry1,carry2,cout;

halfadder_nor HA1 (cout,carry1,r,s);
halfadder_nor HA2 (c0,carry2,cout,t);
or_nor OR1 (c1,carry1,carry2);

endmodule // full_adder




// -------------------------------
// -- half adder with NOR gate
// -------------------------------

module halfadder_nor (s0, s1, a, b);
 output s0,s1;
 input  a, b;
 
  xor_nor XOR1 (s0,a,b);
  and_nor AND1 (s1,a,b);

endmodule // halfadder_nor

// ---------------------
// -- xor with NOR gate
// ---------------------

module xor_nor (s, a, b);
 output s;
 input  a, b;
 wire temp1,temp2,temp3,temp4,temp5,temp6;
 
  nor NOR1 (temp1,b,b);
  nor NOR2 (temp2,a,a);
  nor NOR3 (temp3,a,temp1);
  nor NOR4 (temp4,b,temp2);
  nor NOR5 (temp5, temp3, temp4); 
  nor NOR6 (s, temp5, temp5); 
  
endmodule // xor_nor


// ---------------------
// -- and with NOR gate
// ---------------------

module and_nor (s, a, b);
 output s;
 input  a, b;
 wire temp1,temp2;
 
  nor NOR1 (temp1,a,a);
  nor NOR2 (temp2,b,b);
  nor NOR3 (s, temp1,temp2);

endmodule // and_nor

// ---------------------
// -- or with NOR gate
// ---------------------

module or_nor (s, a, b);
 output s;
 input  a, b;
 wire temp1;
 
  nor NOR1 (temp1,a,b);
  nor NOR2 (s,temp1,temp1);
  
endmodule // or_nor


// -----------------------------
// -- test 4_bits_fulladder_with_nor
// -----------------------------

module test;
 reg [3:0]  a;
 reg [3:0]  b;
 wire [4:0] c;
 integer i,j;
          
// instancia
 four_bits_fulladder_nor FBFA1 (c,a,b);
 
initial begin:start
      a=0; b=0;
 end
 
 
 // parte principal
 initial begin:main
      $display("Guia 05_01 - Alyson Deives - 416589");
      $display("FULL ADDER de 4 bits com portas NOR\n");
		$display("\n   A   +   B  =   S  \n");
		$monitor("  %b%b%b%b + %b%b%b%b = %b%b%b%b%b", a[3],a[2],a[1],a[0],b[3],b[2],b[1],b[0],c[4],c[3],c[2],c[1],c[0]); 
  for(i=0;i<=15;i=i+1) 
  	begin
	
  		for(j=0;j<=15;j=j+1) 
  			begin
			#1 a = i;b=j;
								 			 
  		end	
  end 
end    

endmodule // testhalfadder_nor


	// -----------------------------
	// -- TESTE
	// -----------------------------
	//--Guia 05_01 - Alyson Deives - 416589
	//--FULL ADDER de 4 bits com portas NOR
	//--    A  +    B =   S
    
    // -- 0000 + 0000 = 00000
    // -- 0000 + 0001 = 00001
    // -- 0000 + 0010 = 00010
    // -- 0000 + 0011 = 00011
    // -- 0000 + 0100 = 00100
    // -- 0000 + 0101 = 00101
    // -- 0000 + 0110 = 00110
    // -- 0000 + 0111 = 00111
    // -- 0000 + 1000 = 01000
    // -- 0000 + 1001 = 01001
    // -- 0000 + 1010 = 01010
    // -- 0000 + 1011 = 01011
    // -- 0000 + 1100 = 01100
    // -- 0000 + 1101 = 01101
    // -- 0000 + 1110 = 01110
    // -- 0000 + 1111 = 01111
    // -- 0001 + 0000 = 00001
    // -- 0001 + 0001 = 00010
    // -- 0001 + 0010 = 00011
    // -- 0001 + 0011 = 00100
    // -- 0001 + 0100 = 00101
    // -- 0001 + 0101 = 00110
    // -- 0001 + 0110 = 00111
    // -- 0001 + 0111 = 01000
    // -- 0001 + 1000 = 01001
    // -- 0001 + 1001 = 01010
    // -- 0001 + 1010 = 01011
    // -- 0001 + 1011 = 01100
    // -- 0001 + 1100 = 01101
    // -- 0001 + 1101 = 01110
    // -- 0001 + 1110 = 01111
    // -- 0001 + 1111 = 10000
    // -- 0010 + 0000 = 00010
    // -- 0010 + 0001 = 00011
    // -- 0010 + 0010 = 00100
    // -- 0010 + 0011 = 00101
    // -- 0010 + 0100 = 00110
    // -- 0010 + 0101 = 00111
    // -- 0010 + 0110 = 01000
    // -- 0010 + 0111 = 01001
    // -- 0010 + 1000 = 01010
    // -- 0010 + 1001 = 01011
    // -- 0010 + 1010 = 01100
    // -- 0010 + 1011 = 01101
    // -- 0010 + 1100 = 01110
    // -- 0010 + 1101 = 01111
    // -- 0010 + 1110 = 10000
    // -- 0010 + 1111 = 10001
    // -- 0011 + 0000 = 00011
    // -- 0011 + 0001 = 00100
    // -- 0011 + 0010 = 00101
    // -- 0011 + 0011 = 00110
    // -- 0011 + 0100 = 00111
    // -- 0011 + 0101 = 01000
    // -- 0011 + 0110 = 01001
    // -- 0011 + 0111 = 01010
    // -- 0011 + 1000 = 01011
    // -- 0011 + 1001 = 01100
    // -- 0011 + 1010 = 01101
    // -- 0011 + 1011 = 01110
    // -- 0011 + 1100 = 01111
    // -- 0011 + 1101 = 10000
    // -- 0011 + 1110 = 10001
    // -- 0011 + 1111 = 10010
    // -- 0100 + 0000 = 00100
    // -- 0100 + 0001 = 00101
    // -- 0100 + 0010 = 00110
    // -- 0100 + 0011 = 00111
    // -- 0100 + 0100 = 01000
    // -- 0100 + 0101 = 01001
    // -- 0100 + 0110 = 01010
    // -- 0100 + 0111 = 01011
    // -- 0100 + 1000 = 01100
    // -- 0100 + 1001 = 01101
    // -- 0100 + 1010 = 01110
    // -- 0100 + 1011 = 01111
    // -- 0100 + 1100 = 10000
    // -- 0100 + 1101 = 10001
    // -- 0100 + 1110 = 10010
    // -- 0100 + 1111 = 10011
    // -- 0101 + 0000 = 00101
    // -- 0101 + 0001 = 00110
    // -- 0101 + 0010 = 00111
    // -- 0101 + 0011 = 01000
    // -- 0101 + 0100 = 01001
    // -- 0101 + 0101 = 01010
    // -- 0101 + 0110 = 01011
    // -- 0101 + 0111 = 01100
    // -- 0101 + 1000 = 01101
    // -- 0101 + 1001 = 01110
    // -- 0101 + 1010 = 01111
    // -- 0101 + 1011 = 10000
    // -- 0101 + 1100 = 10001
    // -- 0101 + 1101 = 10010
    // -- 0101 + 1110 = 10011
    // -- 0101 + 1111 = 10100
    // -- 0110 + 0000 = 00110
    // -- 0110 + 0001 = 00111
    // -- 0110 + 0010 = 01000
    // -- 0110 + 0011 = 01001
    // -- 0110 + 0100 = 01010
    // -- 0110 + 0101 = 01011
    // -- 0110 + 0110 = 01100
    // -- 0110 + 0111 = 01101
    // -- 0110 + 1000 = 01110
    // -- 0110 + 1001 = 01111
    // -- 0110 + 1010 = 10000
    // -- 0110 + 1011 = 10001
    // -- 0110 + 1100 = 10010
    // -- 0110 + 1101 = 10011
    // -- 0110 + 1110 = 10100
    // -- 0110 + 1111 = 10101
    // -- 0111 + 0000 = 00111
    // -- 0111 + 0001 = 01000
    // -- 0111 + 0010 = 01001
    // -- 0111 + 0011 = 01010
    // -- 0111 + 0100 = 01011
    // -- 0111 + 0101 = 01100
    // -- 0111 + 0110 = 01101
    // -- 0111 + 0111 = 01110
    // -- 0111 + 1000 = 01111
    // -- 0111 + 1001 = 10000
    // -- 0111 + 1010 = 10001
    // -- 0111 + 1011 = 10010
    // -- 0111 + 1100 = 10011
    // -- 0111 + 1101 = 10100
    // -- 0111 + 1110 = 10101
    // -- 0111 + 1111 = 10110
    // -- 1000 + 0000 = 01000
    // -- 1000 + 0001 = 01001
    // -- 1000 + 0010 = 01010
    // -- 1000 + 0011 = 01011
    // -- 1000 + 0100 = 01100
    // -- 1000 + 0101 = 01101
    // -- 1000 + 0110 = 01110
    // -- 1000 + 0111 = 01111
    // -- 1000 + 1000 = 10000
    // -- 1000 + 1001 = 10001
    // -- 1000 + 1010 = 10010
    // -- 1000 + 1011 = 10011
    // -- 1000 + 1100 = 10100
    // -- 1000 + 1101 = 10101
    // -- 1000 + 1110 = 10110
    // -- 1000 + 1111 = 10111
    // -- 1001 + 0000 = 01001
    // -- 1001 + 0001 = 01010
    // -- 1001 + 0010 = 01011
    // -- 1001 + 0011 = 01100
    // -- 1001 + 0100 = 01101
    // -- 1001 + 0101 = 01110
    // -- 1001 + 0110 = 01111
    // -- 1001 + 0111 = 10000
    // -- 1001 + 1000 = 10001
    // -- 1001 + 1001 = 10010
    // -- 1001 + 1010 = 10011
    // -- 1001 + 1011 = 10100
    // -- 1001 + 1100 = 10101
    // -- 1001 + 1101 = 10110
    // -- 1001 + 1110 = 10111
    // -- 1001 + 1111 = 11000
    // -- 1010 + 0000 = 01010
    // -- 1010 + 0001 = 01011
    // -- 1010 + 0010 = 01100
    // -- 1010 + 0011 = 01101
    // -- 1010 + 0100 = 01110
    // -- 1010 + 0101 = 01111
    // -- 1010 + 0110 = 10000
    // -- 1010 + 0111 = 10001
    // -- 1010 + 1000 = 10010
    // -- 1010 + 1001 = 10011
    // -- 1010 + 1010 = 10100
    // -- 1010 + 1011 = 10101
    // -- 1010 + 1100 = 10110
    // -- 1010 + 1101 = 10111
    // -- 1010 + 1110 = 11000
    // -- 1010 + 1111 = 11001
    // -- 1011 + 0000 = 01011
    // -- 1011 + 0001 = 01100
    // -- 1011 + 0010 = 01101
    // -- 1011 + 0011 = 01110
    // -- 1011 + 0100 = 01111
    // -- 1011 + 0101 = 10000
    // -- 1011 + 0110 = 10001
    // -- 1011 + 0111 = 10010
    // -- 1011 + 1000 = 10011
    // -- 1011 + 1001 = 10100
    // -- 1011 + 1010 = 10101
    // -- 1011 + 1011 = 10110
    // -- 1011 + 1100 = 10111
    // -- 1011 + 1101 = 11000
    // -- 1011 + 1110 = 11001
    // -- 1011 + 1111 = 11010
    // -- 1100 + 0000 = 01100
    // -- 1100 + 0001 = 01101
    // -- 1100 + 0010 = 01110
    // -- 1100 + 0011 = 01111
    // -- 1100 + 0100 = 10000
    // -- 1100 + 0101 = 10001
    // -- 1100 + 0110 = 10010
    // -- 1100 + 0111 = 10011
    // -- 1100 + 1000 = 10100
    // -- 1100 + 1001 = 10101
    // -- 1100 + 1010 = 10110
    // -- 1100 + 1011 = 10111
    // -- 1100 + 1100 = 11000
    // -- 1100 + 1101 = 11001
    // -- 1100 + 1110 = 11010
    // -- 1100 + 1111 = 11011
    // -- 1101 + 0000 = 01101
    // -- 1101 + 0001 = 01110
    // -- 1101 + 0010 = 01111
    // -- 1101 + 0011 = 10000
    // -- 1101 + 0100 = 10001
    // -- 1101 + 0101 = 10010
    // -- 1101 + 0110 = 10011
    // -- 1101 + 0111 = 10100
    // -- 1101 + 1000 = 10101
    // -- 1101 + 1001 = 10110
    // -- 1101 + 1010 = 10111
    // -- 1101 + 1011 = 11000
    // -- 1101 + 1100 = 11001
    // -- 1101 + 1101 = 11010
    // -- 1101 + 1110 = 11011
    // -- 1101 + 1111 = 11100
    // -- 1110 + 0000 = 01110
    // -- 1110 + 0001 = 01111
    // -- 1110 + 0010 = 10000
    // -- 1110 + 0011 = 10001
    // -- 1110 + 0100 = 10010
    // -- 1110 + 0101 = 10011
    // -- 1110 + 0110 = 10100
    // -- 1110 + 0111 = 10101
    // -- 1110 + 1000 = 10110
    // -- 1110 + 1001 = 10111
    // -- 1110 + 1010 = 11000
    // -- 1110 + 1011 = 11001
    // -- 1110 + 1100 = 11010
    // -- 1110 + 1101 = 11011
    // -- 1110 + 1110 = 11100
    // -- 1110 + 1111 = 11101
    // -- 1111 + 0000 = 01111
    // -- 1111 + 0001 = 10000
    // -- 1111 + 0010 = 10001
    // -- 1111 + 0011 = 10010
    // -- 1111 + 0100 = 10011
    // -- 1111 + 0101 = 10100
    // -- 1111 + 0110 = 10101
    // -- 1111 + 0111 = 10110
    // -- 1111 + 1000 = 10111
    // -- 1111 + 1001 = 11000
    // -- 1111 + 1010 = 11001
    // -- 1111 + 1011 = 11010
    // -- 1111 + 1100 = 11011
    // -- 1111 + 1101 = 11100
    // -- 1111 + 1110 = 11101
    // -- 1111 + 1111 = 11110