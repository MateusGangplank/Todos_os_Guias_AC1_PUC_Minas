// Exercicio10 - OR c/ 3 entradas
// Nome: Marlon Henrique de Azeredo Formiga 
// Matricula: 397248 
// ------------------------- 
// ------------------------- 
// -- or gate 
// ------------------------- 

// UMA SAIDA, NAO DUAS !

module orgate ( output s,
						output t,
						input p, 
						input q,
						input r); 
assign s = p | q;
assign t = s | r; 
endmodule // orgate 
// --------------------- 
// -- test or gate 
// --------------------- 
module testorgate; 
// ------------------------- dados locais 
reg a, b, c; // definir registradores 
wire s, t; // definir conexao (fio) 
// ------------------------- instancia 
orgate OR1 (s, t, a, b, c); 
// ------------------------- preparacao 
initial begin:start 
// atribuicao simultanea dos valores iniciais 
a=0; b=0; c=0;
end 
// ------------------------- parte principal 
initial begin 
$display("Exercicio10 - Marlon Henrique de Azeredo Formiga - 397248"); 
$display("Test OR gate"); 
$display("\n(a | b) | c = s\n"); 
a=0; b=0; c=0;
#1 $display("(%b | %b) | %b = %b", a, b, c, t); 
a=1; b=0; c=0;
#1 $display("(%b | %b) | %b = %b", a, b, c, t); 
a=0; b=1; c=0;
#1 $display("(%b | %b) | %b = %b", a, b, c, t);
a=0; b=0; c=1; 
#1 $display("(%b | %b) | %b = %b", a, b, c, t);
a=1; b=1; c=0; 
#1 $display("(%b | %b) | %b = %b", a, b, c, t);
a=0; b=1; c=1;
#1 $display("(%b | %b) | %b = %b", a, b, c, t);
a=1; b=0; c=1;
#1 $display("(%b | %b) | %b = %b", a, b, c, t); 
a=1; b=1; c=1;
#1 $display("(%b | %b) | %b = %b", a, b, c, t); 
end 
endmodule // testorgate 