// --------------------- 
// Exercicio0012 - UM 
// Nome: Marcio Enio G Dutra Junior 
// Matricula: 441698 
// --------------------- 
 
// --------------------- 
// -- um 
// --------------------- 
 
module um (output s, input[7:0] p); 
	assign s = p[0]|p[1]|p[2]|p[3]|p[4]|p[5]|p[6]|p[7]; 
endmodule // um 
 
// --------------------- 
// -- test um
// --------------------- 
module testum; 
// ------------------------- dados locais 
   reg[7:0]   a; // definir registrador 
   wire  s;    // definir conexao (fio) 
// ------------------------- instancia 
   um UM1(s, a);
 
// ------------------------- preparacao 
   initial begin:start 
            a=8'b0000_0000; 
   end 
 
// ------------------------- parte principal 
   initial begin:main 
         $display("Exercicio0012 - Marcio Enio G Dutra Junior - 441698"); 
         $display("Test um"); 
         $display("\np  =  s\n"); 
 	#1    $monitor("%b  =  %b", a, s); 
	#1		a=8'b0000_0001;
	#1		a=8'b0000_0010;
	#1		a=8'b0000_0011;
	#1		a=8'b0000_0100;
	#1		a=8'b0000_0101;
	#1		a=8'b0000_0110;
	#1		a=8'b0000_0111;
	#1		a=8'b0000_1000;
	#1		a=8'b0000_1001;
	#1		a=8'b0000_1010;
	#1		a=8'b0000_1011;
	#1		a=8'b0000_1100;
	#1		a=8'b0000_1101;
	#1		a=8'b0000_1110;
	#1		a=8'b1111_1111;
 
 end 
 
endmodule // testum