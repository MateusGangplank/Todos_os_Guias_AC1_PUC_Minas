Arial// -------------------------
// Exemplo0021 � FULL ADDER
// Nome: Fabio Fiuza Pereira
// Matricula: 406087
// -------------------------
// -------------------------
// full adder
// -------------------------
module fullAdder (output s,
input a,
input b,
input carryIn);
// descrever por portas
endmodule // fullAdder
module test_fullAdder;
// ------------------------- definir dados
reg [2:0] x;
reg [2:0] y;
reg carry;
wire [2:0] soma;
// ------------------------- parte principal
initial begin
$display("Exemplo0021 - xxx yyy zzz - 999999");
$display("Test ALU�s full adder");
// projetar testes do somador complete
end
endmodule // test_fullAdder