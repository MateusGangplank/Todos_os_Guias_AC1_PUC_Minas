// Guia 05
// Nome: Raphaela Fernanda Silva
// Matricula: 420141

module operadorMS ( s4, s3, a, b);
output s4, s3;
input a, b;

xor XOR2(s4,a,b);
and AND2(s3,a,b);

endmodule

module operadorSC ( s0, s1, a, b, v1 );
output s0, s1;
input a, b, v1;
wire s3, s4;

operadorMS MS1(s4,s3,a,b);
operadorMS MS2( s0, s2 ,v1 ,s4);
or OR1(s1,s2,s3);

endmodule

module SC4Bits ( s, a, b);
output[4:0]s;
input[3:0]a,b;
wire[2:0]c;

operadorMS MS1(s[0],c[0],a[0],b[0]);
operadorSC SC1(s[1],c[1],a[1],b[1],c[0]);
operadorSC SC2(s[2],c[2],a[2],b[2],c[1]);
operadorSC SC3(s[3],s[4],a[3],b[3],c[2]);

endmodule


module testSC;
reg [3:0]a,b;
wire [4:0]s;
integer i, j;

SC4Bits SC4B(s, a, b);

 initial begin : start
 
 a=0; b=0;
 
 end

initial begin : main

#1 $display ( " Operador Soma Completa - 4 Bits " );
#1 $display ( "   a  +  b   =  s   " );
	$monitor ( " %4b  %4b  = %5b ",a,b,s);
	
	for ( i = 0; i < 16; i = i + 1)begin
	 a = i;
	for ( j = 0; j < 16; j = j + 1)begin
	#1 b = j;
	end
	end
				
end

endmodule

/* Operador Soma Completa - 4 Bits 
       a  +  b   =  s   
     0000  0000  = 00000 
     0000  0001  = 00001 
     0000  0010  = 00010 
     0000  0011  = 00011 
     0000  0100  = 00100 
     0000  0101  = 00101 
     0000  0110  = 00110 
     0000  0111  = 00111 
     0000  1000  = 01000 
     0000  1001  = 01001 
     0000  1010  = 01010 
     0000  1011  = 01011 
     0000  1100  = 01100 
     0000  1101  = 01101 
     0000  1110  = 01110 
     0001  1111  = 10000 
     0001  0000  = 00001 
     0001  0001  = 00010 
     0001  0010  = 00011 
     0001  0011  = 00100 
     0001  0100  = 00101 
     0001  0101  = 00110 
     0001  0110  = 00111 
     0001  0111  = 01000 
     0001  1000  = 01001 
     0001  1001  = 01010 
     0001  1010  = 01011 
     0001  1011  = 01100 
     0001  1100  = 01101 
     0001  1101  = 01110 
     0001  1110  = 01111 
     0010  1111  = 10001 
     0010  0000  = 00010 
     0010  0001  = 00011 
     0010  0010  = 00100 
     0010  0011  = 00101 
     0010  0100  = 00110 
     0010  0101  = 00111 
     0010  0110  = 01000 
     0010  0111  = 01001 
     0010  1000  = 01010 
     0010  1001  = 01011 
     0010  1010  = 01100 
     0010  1011  = 01101 
     0010  1100  = 01110 
     0010  1101  = 01111 
     0010  1110  = 10000 
     0011  1111  = 10010 
     0011  0000  = 00011 
     0011  0001  = 00100 
     0011  0010  = 00101 
     0011  0011  = 00110 
     0011  0100  = 00111 
     0011  0101  = 01000 
     0011  0110  = 01001 
     0011  0111  = 01010 
     0011  1000  = 01011 
     0011  1001  = 01100 
     0011  1010  = 01101 
     0011  1011  = 01110 
     0011  1100  = 01111 
     0011  1101  = 10000 
     0011  1110  = 10001 
     0100  1111  = 10011 
     0100  0000  = 00100 
     0100  0001  = 00101 
     0100  0010  = 00110 
     0100  0011  = 00111 
     0100  0100  = 01000 
     0100  0101  = 01001 
     0100  0110  = 01010 
     0100  0111  = 01011 
     0100  1000  = 01100 
     0100  1001  = 01101 
     0100  1010  = 01110 
     0100  1011  = 01111 
     0100  1100  = 10000 
     0100  1101  = 10001 
     0100  1110  = 10010 
     0101  1111  = 10100 
     0101  0000  = 00101 
     0101  0001  = 00110 
     0101  0010  = 00111 
     0101  0011  = 01000 
     0101  0100  = 01001 
     0101  0101  = 01010 
     0101  0110  = 01011 
     0101  0111  = 01100 
     0101  1000  = 01101 
     0101  1001  = 01110 
     0101  1010  = 01111 
     0101  1011  = 10000 
     0101  1100  = 10001 
     0101  1101  = 10010 
     0101  1110  = 10011 
     0110  1111  = 10101 
     0110  0000  = 00110 
     0110  0001  = 00111 
     0110  0010  = 01000 
     0110  0011  = 01001 
     0110  0100  = 01010 
     0110  0101  = 01011 
     0110  0110  = 01100 
     0110  0111  = 01101 
     0110  1000  = 01110 
     0110  1001  = 01111 
     0110  1010  = 10000 
     0110  1011  = 10001 
     0110  1100  = 10010 
     0110  1101  = 10011 
     0110  1110  = 10100 
     0111  1111  = 10110 
     0111  0000  = 00111 
     0111  0001  = 01000 
     0111  0010  = 01001 
     0111  0011  = 01010 
     0111  0100  = 01011 
     0111  0101  = 01100 
     0111  0110  = 01101 
     0111  0111  = 01110 
     0111  1000  = 01111 
     0111  1001  = 10000 
     0111  1010  = 10001 
     0111  1011  = 10010 
     0111  1100  = 10011 
     0111  1101  = 10100 
     0111  1110  = 10101 
     1000  1111  = 10111 
     1000  0000  = 01000 
     1000  0001  = 01001 
     1000  0010  = 01010 
     1000  0011  = 01011 
     1000  0100  = 01100 
     1000  0101  = 01101 
     1000  0110  = 01110 
     1000  0111  = 01111 
     1000  1000  = 10000 
     1000  1001  = 10001 
     1000  1010  = 10010 
     1000  1011  = 10011 
     1000  1100  = 10100 
     1000  1101  = 10101 
     1000  1110  = 10110 
     1001  1111  = 11000 
     1001  0000  = 01001 
     1001  0001  = 01010 
     1001  0010  = 01011 
     1001  0011  = 01100 
     1001  0100  = 01101 
     1001  0101  = 01110 
     1001  0110  = 01111 
     1001  0111  = 10000 
     1001  1000  = 10001 
     1001  1001  = 10010 
     1001  1010  = 10011 
     1001  1011  = 10100 
     1001  1100  = 10101 
     1001  1101  = 10110 
     1001  1110  = 10111 
     1010  1111  = 11001 
     1010  0000  = 01010 
     1010  0001  = 01011 
     1010  0010  = 01100 
     1010  0011  = 01101 
     1010  0100  = 01110 
     1010  0101  = 01111 
     1010  0110  = 10000 
     1010  0111  = 10001 
     1010  1000  = 10010 
     1010  1001  = 10011 
     1010  1010  = 10100 
     1010  1011  = 10101 
     1010  1100  = 10110 
     1010  1101  = 10111 
    
     1010  1110  = 11000 
     1011  1111  = 11010 
     1011  0000  = 01011 
     1011  0001  = 01100 
     1011  0010  = 01101 
     1011  0011  = 01110 
     1011  0100  = 01111 
     1011  0101  = 10000 
     1011  0110  = 10001 
     1011  0111  = 10010 
     1011  1000  = 10011 
     1011  1001  = 10100 
     1011  1010  = 10101 
     1011  1011  = 10110 
     1011  1100  = 10111 
     1011  1101  = 11000 
     1011  1110  = 11001 
     1100  1111  = 11011 
     1100  0000  = 01100 
     1100  0001  = 01101 
     1100  0010  = 01110 
     1100  0011  = 01111 
     1100  0100  = 10000 
     1100  0101  = 10001 
     1100  0110  = 10010 
     1100  0111  = 10011 
     1100  1000  = 10100 
     1100  1001  = 10101 
     1100  1010  = 10110 
     1100  1011  = 10111 
     1100  1100  = 11000 
     1100  1101  = 11001 
     1100  1110  = 11010 
     1101  1111  = 11100 
     1101  0000  = 01101 
     1101  0001  = 01110 
     1101  0010  = 01111 
     1101  0011  = 10000 
     1101  0100  = 10001 
     1101  0101  = 10010 
     1101  0110  = 10011 
     1101  0111  = 10100 
     1101  1000  = 10101 
     1101  1001  = 10110 
     1101  1010  = 10111 
     1101  1011  = 11000 
     1101  1100  = 11001 
     1101  1101  = 11010 
     1101  1110  = 11011 
     1110  1111  = 11101 
     1110  0000  = 01110 
     1110  0001  = 01111 
     1110  0010  = 10000 
     1110  0011  = 10001 
     1110  0100  = 10010 
     1110  0101  = 10011 
     1110  0110  = 10100 
     1110  0111  = 10101 
     1110  1000  = 10110 
     1110  1001  = 10111 
     1110  1010  = 11000 
     1110  1011  = 11001 
     1110  1100  = 11010 
     1110  1101  = 11011 
     1110  1110  = 11100 
     1111  1111  = 11110 
     1111  0000  = 01111 
     1111  0001  = 10000 
     1111  0010  = 10001 
     1111  0011  = 10010 
     1111  0100  = 10011 
     1111  0101  = 10100 
     1111  0110  = 10101 
     1111  0111  = 10110 
     1111  1000  = 10111 
     1111  1001  = 11000 
     1111  1010  = 11001 
     1111  1011  = 11010 
     1111  1100  = 11011 
     1111  1101  = 11100 
     1111  1110  = 11101 
     1111  1111  = 11110 
*/
