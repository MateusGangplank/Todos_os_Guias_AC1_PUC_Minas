//Nome: Vitor Angelo Lima
//Matricula: 451621
module clock ( clk );
	output clk;
	reg clk;
	initial begin
		clk = 1'b0;
	end

	always begin
		#1 clk = ~clk;
	end
endmodule // clock ( )
