// ------------------------- 
// Guia08_04 - Registrador de Deslocamento
// Nome: Bruno Cezar Andrade Viallet 
// Matricula: 396679
// ------------------------- 


//-----------------------------
// -- CLOCK
//-----------------------------
`include "clock.v"


// -------------------------
// -- FLIP FLOP D
// -------------------------
module ffd(q,qnot,data,clk);
	output q;
	output qnot;
	input data;
	input clk;
	
	reg q,qnot;
	
	initial begin
		q = 1'b0;
		qnot = 1'b1;
	end
	always @ (posedge clk)
		begin
		q <= data;	qnot <= ~q;
		end
			
endmodule //ffd

// --------------------------------------------------------------------------------------------------
// --  Registrador de deslocamento circular, em anel torcido, para a esquerda, 4bits
// --------------------------------------------------------------------------------------------------
module rotateLeftRegister (output [3:0]s, input d, input clk);
wire nots;	
	
	or OR1 (d0, d, s[3]);
	
	ffd FF0 (s[0], nots, d0, clk);
	ffd FF1 (s[1], nots, s[0], clk);
	ffd FF2 (s[2], nots, s[1], clk);
	ffd FF3 (s[3], nots, s[2], clk);

	
endmodule//rotateLeftRegister

// -------------------------
// -- Teste
// -------------------------

module teste;
wire [3:0] saida;
reg d;
wire clock; 
clock clk ( clock ); 
rotateLeftRegister RLF1 (saida, d, clock);
	
	initial begin
		$display("Guia08_04 - Bruno Cezar Andrade Viallet - 396679"); 
		$display("D CLOCK SAIDA");
		d = 1;
		$monitor("%1b    %1b    %5b", d, clock, saida);
		#23 d = 0;
		#240 $finish;
	end

endmodule //teste
