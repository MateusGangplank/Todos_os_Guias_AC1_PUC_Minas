// ---------------------------
// Guia 09
// ---------------------------

`include "clock.v"

module pulse1 ( signal, clock );
 input  clock;
 output signal;
 reg    signal;

 always @ ( negedge clock )
  begin
      signal = 1'b1;
  #60  signal = 1'b0;
  end
endmodule // pulse

module Guia0904;

 wire  clock;
 clock clk ( clock );
 wire  p1;

 pulse1   pls1   ( p1, clock );

 initial begin
  $dumpfile ( "Guia0904.vcd" );
  $dumpvars ( 1, clock, p1);

  #480 $finish;
 end

endmodule
