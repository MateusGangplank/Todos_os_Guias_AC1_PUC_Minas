// ---------------------
// Guia 05_01 - Soma Completa 4 bits
// Nome: Anderson Belchior de Carvalho
// Matricula: 396673
// ---------------------

// ---------------------
// -- meia soma
// ---------------------

module meiasoma (s, v, p, q);

output v, s;
input p, q;

xor XOR1 (s, p, q);
and AND1 (v, p, q);

endmodule // meisoma

// ---------------------
// -- soma completa
// ---------------------

module somacompleta (s0, s1, p, q, v);

output s1, s0;
input p, q, v;
wire t1, t2, t3;

MS MS1 (t2, t1, p, q);
MS MS2 (s0, t3, v, t2);
or Or1 (s1, t3, t1);

endmodule // somacompleta


module metodoSomador4bits(saida,carryout,e1,e2);

output [3:0]saida;
output carryout;
input [3:0]e1,e2;
wire carryout1,carryout2,carryout3;

metodomeiasoma MEIASOMA (saida[0],carryout1,e1[0],e2[0]);
metodosomacompleta SOMACOMPLETA1 (saida[1],carryout2,e1[1],e2[1],carryout1);
metodosomacompleta SOMACOMPLETA2 (saida[2],carryout3,e1[2],e2[2],carryout2);
metodosomacompleta SOMACOMPLETA3 (saida[3],carryout,e1[3],e2[3],carryout3);

endmodule


module testsomador4bits;
reg [3:0]e1,e2;
wire [3:0]saida;
wire carry;
integer i,j;

metodoSomador4bits Somador4bits(saida,carry,e1,e2);

initial begin: start
		e1=0; e2=0;
end


	initial begin:main

		$display("Circuito Soma Completa com 4 bits ");
		#1 $display(" e1 + e2 = carry saida ");
		#1 $monitor(" %4b + %4b = %b %4b", e1,e2,carry,saida);

		for( i=0; i<=15; i = i+1 )
		begin
			e1 = i;
			for ( j=0; j<=15; j = j+1 )
			begin
				#1 e2 = j;
			end
		end

	end

endmodule

/* Registrando os resultados

  
    Circuito Soma Completa com 4 bits 
     e1 + e2 = carry saida 
     0000 + 0000 = 0 0000
     0000 + 0001 = 0 0001
     0000 + 0010 = 0 0010
     0000 + 0011 = 0 0011
     0000 + 0100 = 0 0100
     0000 + 0101 = 0 0101
     0000 + 0110 = 0 0110
     0000 + 0111 = 0 0111
     0000 + 1000 = 0 1000
     0000 + 1001 = 0 1001
     0000 + 1010 = 0 1010
     0000 + 1011 = 0 1011
     0000 + 1100 = 0 1100
     0000 + 1101 = 0 1101
     0000 + 1110 = 0 1110
     0001 + 1111 = 1 0000
     0001 + 0000 = 0 0001
     0001 + 0001 = 0 0010
     0001 + 0010 = 0 0011
     0001 + 0011 = 0 0100
     0001 + 0100 = 0 0101
     0001 + 0101 = 0 0110
     0001 + 0110 = 0 0111
     0001 + 0111 = 0 1000
     0001 + 1000 = 0 1001
     0001 + 1001 = 0 1010
     0001 + 1010 = 0 1011
     0001 + 1011 = 0 1100
     0001 + 1100 = 0 1101
     0001 + 1101 = 0 1110
     0001 + 1110 = 0 1111
     0010 + 1111 = 1 0001
     0010 + 0000 = 0 0010
     0010 + 0001 = 0 0011
     0010 + 0010 = 0 0100
     0010 + 0011 = 0 0101
     0010 + 0100 = 0 0110
     0010 + 0101 = 0 0111
     0010 + 0110 = 0 1000
     0010 + 0111 = 0 1001
     0010 + 1000 = 0 1010
     0010 + 1001 = 0 1011
     0010 + 1010 = 0 1100
     0010 + 1011 = 0 1101
     0010 + 1100 = 0 1110
     0010 + 1101 = 0 1111
     0010 + 1110 = 1 0000
     0011 + 1111 = 1 0010
     0011 + 0000 = 0 0011
     0011 + 0001 = 0 0100
     0011 + 0010 = 0 0101
     0011 + 0011 = 0 0110
     0011 + 0100 = 0 0111
     0011 + 0101 = 0 1000
     0011 + 0110 = 0 1001
     0011 + 0111 = 0 1010
     0011 + 1000 = 0 1011
     0011 + 1001 = 0 1100
     0011 + 1010 = 0 1101
     0011 + 1011 = 0 1110
     0011 + 1100 = 0 1111
     0011 + 1101 = 1 0000
     0011 + 1110 = 1 0001
     0100 + 1111 = 1 0011
     0100 + 0000 = 0 0100
     0100 + 0001 = 0 0101
     0100 + 0010 = 0 0110
     0100 + 0011 = 0 0111
     0100 + 0100 = 0 1000
     0100 + 0101 = 0 1001
     0100 + 0110 = 0 1010
     0100 + 0111 = 0 1011
     0100 + 1000 = 0 1100
     0100 + 1001 = 0 1101
     0100 + 1010 = 0 1110
     0100 + 1011 = 0 1111
     0100 + 1100 = 1 0000
     0100 + 1101 = 1 0001
     0100 + 1110 = 1 0010
     0101 + 1111 = 1 0100
     0101 + 0000 = 0 0101
     0101 + 0001 = 0 0110
     0101 + 0010 = 0 0111
     0101 + 0011 = 0 1000
     0101 + 0100 = 0 1001
     0101 + 0101 = 0 1010
     0101 + 0110 = 0 1011
     0101 + 0111 = 0 1100
     0101 + 1000 = 0 1101
     0101 + 1001 = 0 1110
     0101 + 1010 = 0 1111
     0101 + 1011 = 1 0000
     0101 + 1100 = 1 0001
     0101 + 1101 = 1 0010
     0101 + 1110 = 1 0011
     0110 + 1111 = 1 0101
     0110 + 0000 = 0 0110
     0110 + 0001 = 0 0111
     0110 + 0010 = 0 1000
     0110 + 0011 = 0 1001
     0110 + 0100 = 0 1010
     0110 + 0101 = 0 1011
     0110 + 0110 = 0 1100
     0110 + 0111 = 0 1101
     0110 + 1000 = 0 1110
     0110 + 1001 = 0 1111
     0110 + 1010 = 1 0000
     0110 + 1011 = 1 0001
     0110 + 1100 = 1 0010
     0110 + 1101 = 1 0011
     0110 + 1110 = 1 0100
     0111 + 1111 = 1 0110
     0111 + 0000 = 0 0111
     0111 + 0001 = 0 1000
     0111 + 0010 = 0 1001
     0111 + 0011 = 0 1010
     0111 + 0100 = 0 1011
     0111 + 0101 = 0 1100
     0111 + 0110 = 0 1101
     0111 + 0111 = 0 1110
     0111 + 1000 = 0 1111
     0111 + 1001 = 1 0000
     0111 + 1010 = 1 0001
     0111 + 1011 = 1 0010
     0111 + 1100 = 1 0011
     0111 + 1101 = 1 0100
     0111 + 1110 = 1 0101
     1000 + 1111 = 1 0111
     1000 + 0000 = 0 1000
     1000 + 0001 = 0 1001
     1000 + 0010 = 0 1010
     1000 + 0011 = 0 1011
     1000 + 0100 = 0 1100
     1000 + 0101 = 0 1101
     1000 + 0110 = 0 1110
     1000 + 0111 = 0 1111
     1000 + 1000 = 1 0000
     1000 + 1001 = 1 0001
     1000 + 1010 = 1 0010
     1000 + 1011 = 1 0011
     1000 + 1100 = 1 0100
     1000 + 1101 = 1 0101
     1000 + 1110 = 1 0110
     1001 + 1111 = 1 1000
     1001 + 0000 = 0 1001
     1001 + 0001 = 0 1010
     1001 + 0010 = 0 1011
     1001 + 0011 = 0 1100
     1001 + 0100 = 0 1101
     1001 + 0101 = 0 1110
     1001 + 0110 = 0 1111
     1001 + 0111 = 1 0000
     1001 + 1000 = 1 0001
     1001 + 1001 = 1 0010
     1001 + 1010 = 1 0011
     1001 + 1011 = 1 0100
     1001 + 1100 = 1 0101
     1001 + 1101 = 1 0110
     1001 + 1110 = 1 0111
     1010 + 1111 = 1 1001
     1010 + 0000 = 0 1010
     1010 + 0001 = 0 1011
     1010 + 0010 = 0 1100
     1010 + 0011 = 0 1101
     1010 + 0100 = 0 1110
     1010 + 0101 = 0 1111
     1010 + 0110 = 1 0000
     1010 + 0111 = 1 0001
     1010 + 1000 = 1 0010
     1010 + 1001 = 1 0011
     1010 + 1010 = 1 0100
     1010 + 1011 = 1 0101
     1010 + 1100 = 1 0110
     1010 + 1101 = 1 0111
    
     1010 + 1110 = 1 1000
     1011 + 1111 = 1 1010
     1011 + 0000 = 0 1011
     1011 + 0001 = 0 1100
     1011 + 0010 = 0 1101
     1011 + 0011 = 0 1110
     1011 + 0100 = 0 1111
     1011 + 0101 = 1 0000
     1011 + 0110 = 1 0001
     1011 + 0111 = 1 0010
     1011 + 1000 = 1 0011
     1011 + 1001 = 1 0100
     1011 + 1010 = 1 0101
     1011 + 1011 = 1 0110
     1011 + 1100 = 1 0111
     1011 + 1101 = 1 1000
     1011 + 1110 = 1 1001
     1100 + 1111 = 1 1011
     1100 + 0000 = 0 1100
     1100 + 0001 = 0 1101
     1100 + 0010 = 0 1110
     1100 + 0011 = 0 1111
     1100 + 0100 = 1 0000
     1100 + 0101 = 1 0001
     1100 + 0110 = 1 0010
     1100 + 0111 = 1 0011
     1100 + 1000 = 1 0100
     1100 + 1001 = 1 0101
     1100 + 1010 = 1 0110
     1100 + 1011 = 1 0111
     1100 + 1100 = 1 1000
     1100 + 1101 = 1 1001
     1100 + 1110 = 1 1010
     1101 + 1111 = 1 1100
     1101 + 0000 = 0 1101
     1101 + 0001 = 0 1110
     1101 + 0010 = 0 1111
     1101 + 0011 = 1 0000
     1101 + 0100 = 1 0001
     1101 + 0101 = 1 0010
     1101 + 0110 = 1 0011
     1101 + 0111 = 1 0100
     1101 + 1000 = 1 0101
     1101 + 1001 = 1 0110
     1101 + 1010 = 1 0111
     1101 + 1011 = 1 1000
     1101 + 1100 = 1 1001
     1101 + 1101 = 1 1010
     1101 + 1110 = 1 1011
     1110 + 1111 = 1 1101
     1110 + 0000 = 0 1110
     1110 + 0001 = 0 1111
     1110 + 0010 = 1 0000
     1110 + 0011 = 1 0001
     1110 + 0100 = 1 0010
     1110 + 0101 = 1 0011
     1110 + 0110 = 1 0100
     1110 + 0111 = 1 0101
     1110 + 1000 = 1 0110
     1110 + 1001 = 1 0111
     1110 + 1010 = 1 1000
     1110 + 1011 = 1 1001
     1110 + 1100 = 1 1010
     1110 + 1101 = 1 1011
     1110 + 1110 = 1 1100
     1111 + 1111 = 1 1110
     1111 + 0000 = 0 1111
     1111 + 0001 = 1 0000
     1111 + 0010 = 1 0001
     1111 + 0011 = 1 0010
     1111 + 0100 = 1 0011
     1111 + 0101 = 1 0100
     1111 + 0110 = 1 0101
     1111 + 0111 = 1 0110
     1111 + 1000 = 1 0111
     1111 + 1001 = 1 1000
     1111 + 1010 = 1 1001
     1111 + 1011 = 1 1010
     1111 + 1100 = 1 1011
     1111 + 1101 = 1 1100
     1111 + 1110 = 1 1101
     1111 + 1111 = 1 1110
    
     ----jGRASP: operation complete.
    
*/

