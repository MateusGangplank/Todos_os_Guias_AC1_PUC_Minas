// Exemplo 01
// Nome: Bruno Rafael Nicolletti
// Matricula: 380752

module circuito (s0, s1, s2, s3, s4, a4, a3, a2, a1, a0);
 output s0, s1, s2, s3, s4;
 input a4, a3, a2, a1, a0;
 
 not NOT1 (s0, a0);
 not NOT2 (s1, a1);
 not NOT3 (s2, a2);
 not NOT4 (s3, a3);
 not NOT5 (s4, a4);
 
endmodule

module testcircuito;
 reg a4, a3, a2, a1, a0;
 wire s0, s1, s2, s3, s4;
 
 circuito CIRC1 (s0, s1, s2, s3, s4, a4, a3, a2, a1, a0);
 
 initial begin
      $display("Exemplo 01 - Bruno Rafael Nicolletti - 380752");
      $display("Test Circuito Complemento de 1");
      $display("\na4 a3 a2 a1 a0 = s4 s3 s2 s1 s0");
		$monitor(" %b  %b  %b  %b  %b =  %b  %b  %b  %b  %b", a4, a3, a2, a1, a0, s4, s3, s2, s1, s0);
	#1 a4=0; a3=0; a2=0; a1=0; a0=0;
	#1 a4=0; a3=0; a2=0; a1=0; a0=1;
	#1 a4=0; a3=0; a2=0; a1=1; a0=0;
	#1 a4=0; a3=0; a2=0; a1=1; a0=1;
	#1 a4=0; a3=0; a2=1; a1=0; a0=0;
	#1 a4=0; a3=0; a2=1; a1=0; a0=1;
	#1 a4=0; a3=0; a2=1; a1=1; a0=0;
	#1 a4=0; a3=0; a2=1; a1=1; a0=1;
	#1 a4=0; a3=1; a2=0; a1=0; a0=0;
	#1 a4=0; a3=1; a2=0; a1=0; a0=1;
	#1 a4=0; a3=1; a2=0; a1=1; a0=0;
	#1 a4=0; a3=1; a2=0; a1=1; a0=1;
	#1 a4=0; a3=1; a2=1; a1=0; a0=0;
	#1 a4=0; a3=1; a2=1; a1=0; a0=1;
	#1 a4=0; a3=1; a2=1; a1=1; a0=0;
	#1 a4=0; a3=1; a2=1; a1=1; a0=1;
	#1 a4=1; a3=0; a2=0; a1=0; a0=0;
	#1 a4=1; a3=0; a2=0; a1=0; a0=1;
	#1 a4=1; a3=0; a2=0; a1=1; a0=0;
	#1 a4=1; a3=0; a2=0; a1=1; a0=1;
	#1 a4=1; a3=0; a2=1; a1=0; a0=0;
	#1 a4=1; a3=0; a2=1; a1=0; a0=1;
	#1 a4=1; a3=0; a2=1; a1=1; a0=0;
	#1 a4=1; a3=0; a2=1; a1=1; a0=1;
	#1 a4=1; a3=1; a2=0; a1=0; a0=0;
	#1 a4=1; a3=1; a2=0; a1=0; a0=1;
	#1 a4=1; a3=1; a2=0; a1=1; a0=0;
	#1 a4=1; a3=1; a2=0; a1=1; a0=1;
	#1 a4=1; a3=1; a2=1; a1=0; a0=0;
	#1 a4=1; a3=1; a2=1; a1=0; a0=1;
	#1 a4=1; a3=1; a2=1; a1=1; a0=0;
	#1 a4=1; a3=1; a2=1; a1=1; a0=1;
	
 end
 
endmodule

//  a4 a3 a2 a1 a0 = s4 s3 s2 s1 s0
     x  x  x  x  x =  x  x  x  x  x
     0  0  0  0  0 =  1  1  1  1  1
     0  0  0  0  1 =  1  1  1  1  0
     0  0  0  1  0 =  1  1  1  0  1
     0  0  0  1  1 =  1  1  1  0  0
     0  0  1  0  0 =  1  1  0  1  1
     0  0  1  0  1 =  1  1  0  1  0
     0  0  1  1  0 =  1  1  0  0  1
     0  0  1  1  1 =  1  1  0  0  0
     0  1  0  0  0 =  1  0  1  1  1
     0  1  0  0  1 =  1  0  1  1  0
     0  1  0  1  0 =  1  0  1  0  1
     0  1  0  1  1 =  1  0  1  0  0
     0  1  1  0  0 =  1  0  0  1  1
     0  1  1  0  1 =  1  0  0  1  0
     0  1  1  1  0 =  1  0  0  0  1
     0  1  1  1  1 =  1  0  0  0  0
     1  0  0  0  0 =  0  1  1  1  1
     1  0  0  0  1 =  0  1  1  1  0
     1  0  0  1  0 =  0  1  1  0  1
     1  0  0  1  1 =  0  1  1  0  0
     1  0  1  0  0 =  0  1  0  1  1
     1  0  1  0  1 =  0  1  0  1  0
     1  0  1  1  0 =  0  1  0  0  1
     1  0  1  1  1 =  0  1  0  0  0
     1  1  0  0  0 =  0  0  1  1  1
     1  1  0  0  1 =  0  0  1  1  0
     1  1  0  1  0 =  0  0  1  0  1
     1  1  0  1  1 =  0  0  1  0  0
     1  1  1  0  0 =  0  0  0  1  1
     1  1  1  0  1 =  0  0  0  1  0
     1  1  1  1  0 =  0  0  0  0  1
     1  1  1  1  1 =  0  0  0  0  0