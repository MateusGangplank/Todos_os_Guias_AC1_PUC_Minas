// ------------------------- 
// Mealy FSM 
// Nome: Lucas Siqueira Chagas 
// Matricula: 380783
// -------------------------

// -------------------- 
// --- Mealy FSM 
// -------------------- 

  `include "Mealy000_111.v" 
 
  module Exemplo0056; 
   reg clk, reset, x; 
   wire m1; 

   mealy000_111 mealy1 ( m1, x, clk, reset ); 

  initial 
   begin 
    $display ( "Time  X  Mealy " );
	  
// initial values 
   clk = 1; 
   reset = 0; 
   x = 0; 

// input signal changing  
   #5 reset = 1; 
   #5 x = 0; //faz
   #5  
   #5 x = 1; //faz
   #5  
   #5 x = 0; //faz
   #5 
   #5 x = 0; //faz
   #5 
	#5 x = 0; //faz
   #5 
   #5 x = 1; //faz

	#30 $finish; 
   end // initial 

always 
   #5 clk = ~clk; 

always @( posedge clk ) 
 begin 
  $display ( "%4d %4b %4b", $time, x, m1); 
end // always at positive edge clocking changing 

endmodule // Exemplo0056
