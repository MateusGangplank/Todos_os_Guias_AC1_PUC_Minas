// -------------------------
// Nome: Marcio Enio Gon�alves Dutra Junior
// Matricula: 441698
// -------------------------

// -------------- 
// --- Mealy FSM 
// -------------- 
 
/* 
                        Mealy FSM Diagram 
                      __________________ 
                     /                    \ 
              1    v   1           0     1 | // found 
   [start] ---> [id1] ---> [id11] ---> [id110] 
     ^  \0      0 |       1 /  ^         0 | // not found 
      \_/        /          \__/         | 
       \________/                      / 
        \                            / 
         \_________________________/ 
*/ 
// constant definitions 
`define found 1 
`define notfound 0 
 
// FSM by Mealy 
module mealy1100 ( y, x, clk, reset ); 
 output y; 
 input   x; 
 input   clk; 
 input   reset; 
 
 reg      y; 
 
 parameter         // state identifiers  
   start    = 3'b000, 
   id1      = 3'b001, 
   id11    = 3'b011, 
   id110  = 3'b010,
	id1100 = 3'b110;
 
   reg [2:0] E1; // current state variables 
   reg [2:0] E2; // next state logic output 
 
 
// next state logic 
   always @( x or E1 ) 
    begin 
     y = `notfound; 
     case ( E1 ) 
      start: 
        if ( x ) 
         E2 = id1; 
        else 
         E2 = start; 
      id1: 
        if ( x ) 
         E2 = id11; 
        else 
         E2 = start; 
      id11: 
        if ( x ) 
         E2 = id11; 
        else 
         E2 = id110; 
      id110: 
        if ( x ) 
         begin 
           E2 =  id1; 
           y  = `notfound; 
         end 
        else 
         begin 
           E2 =  id1100; 
           y  = `found; 
         end 
		id1100:
			if ( x ) 
         begin 
           E2 =  id1100; 
           y  = `notfound; 
         end 
        else 
         begin 
           E2 =  id1100; 
           y  = `notfound; 
         end 
      default:   // undefined state 
           E2 =  3'bxxx; 
     endcase 
    end // always at signal or state changing 
 
// state variables 
   always @( posedge clk or negedge reset ) 
    begin 
     if ( reset ) 
      E1 = E2;    // updates current state 
     else 
      E1 = 0;     // reset 
    end // always at signal changing 
 
endmodule // mealy1101