// ------------------------------------
// Exemplo0044 - DIFEREN�A
// Nome:Mateus Guilherme do Carmo Cruz
// Matricula: 427446
// ------------------------------------


module funcao(output s, input[3:0]x, input[3:0]y);
	wire [3:0]aux;
	xnor xnor1(aux[0],x[0],y[0]);
	xnor xnor2(aux[1],x[1],y[1]);
	xnor xnor3(aux[2],x[2],y[2]);
	xnor xnor4(aux[3],x[3],y[3]);
	nand nand1(s,aux[0],aux[1],aux[2],aux[3]);
endmodule //funcao

module principal;
	reg [3:0]a,b;
	wire s;
	
	funcao f1(s,a,b);
	
	initial begin
		a = 0; b = 0;
		$display("Exemplo0044 - Mateus Guilherme do Carmo Cruz - 427446"); 
		$display("Test LU's different");
		$display("  a  -   b  =    s");
		$monitor("%4b - %4b = %4b",a,b,s);
		#1 b = 1; #1 b = 2; #1 b = 3; #1 b = 4;
		#1 b = 5; #1 b = 6; #1 b = 7; #1 b = 8;
		#1 b = 9; #1 b = 10; #1 b = 11; #1 b = 12;
		#1 b = 13; #1 b = 14; #1 b = 15;
		
		#1 a = 1; b = 0;
		#1 b = 1; #1 b = 2; #1 b = 3; #1 b = 4;
		#1 b = 5; #1 b = 6; #1 b = 7; #1 b = 8;
		#1 b = 9; #1 b = 10; #1 b = 11; #1 b = 12;
		#1 b = 13; #1 b = 14; #1 b = 15;
		
		#1 a = 2; b = 0;
		#1 b = 1; #1 b = 2; #1 b = 3; #1 b = 4;
		#1 b = 5; #1 b = 6; #1 b = 7; #1 b = 8;
		#1 b = 9; #1 b = 10; #1 b = 11; #1 b = 12;
		#1 b = 13; #1 b = 14; #1 b = 15;
		
		#1 a = 3; b = 0;
		#1 b = 1; #1 b = 2; #1 b = 3; #1 b = 4;
		#1 b = 5; #1 b = 6; #1 b = 7; #1 b = 8;
		#1 b = 9; #1 b = 10; #1 b = 11; #1 b = 12;
		#1 b = 13; #1 b = 14; #1 b = 15;
		
		#1 a = 4; b = 0;
		#1 b = 1; #1 b = 2; #1 b = 3; #1 b = 4;
		#1 b = 5; #1 b = 6; #1 b = 7; #1 b = 8;
		#1 b = 9; #1 b = 10; #1 b = 11; #1 b = 12;
		#1 b = 13; #1 b = 14; #1 b = 15;
		
		#1 a = 5; b = 0;
		#1 b = 1; #1 b = 2; #1 b = 3; #1 b = 4;
		#1 b = 5; #1 b = 6; #1 b = 7; #1 b = 8;
		#1 b = 9; #1 b = 10; #1 b = 11; #1 b = 12;
		#1 b = 13; #1 b = 14; #1 b = 15;
		
		#1 a = 6; b = 0;
		#1 b = 1; #1 b = 2; #1 b = 3; #1 b = 4;
		#1 b = 5; #1 b = 6; #1 b = 7; #1 b = 8;
		#1 b = 9; #1 b = 10; #1 b = 11; #1 b = 12;
		#1 b = 13; #1 b = 14; #1 b = 15;
		
		#1 a = 7; b = 0;
		#1 b = 1; #1 b = 2; #1 b = 3; #1 b = 4;
		#1 b = 5; #1 b = 6; #1 b = 7; #1 b = 8;
		#1 b = 9; #1 b = 10; #1 b = 11; #1 b = 12;
		#1 b = 13; #1 b = 14; #1 b = 15;
		
		#1 a = 8; b = 0;
		#1 b = 1; #1 b = 2; #1 b = 3; #1 b = 4;
		#1 b = 5; #1 b = 6; #1 b = 7; #1 b = 8;
		#1 b = 9; #1 b = 10; #1 b = 11; #1 b = 12;
		#1 b = 13; #1 b = 14; #1 b = 15;
		
		#1 a = 9; b = 0;
		#1 b = 1; #1 b = 2; #1 b = 3; #1 b = 4;
		#1 b = 5; #1 b = 6; #1 b = 7; #1 b = 8;
		#1 b = 9; #1 b = 10; #1 b = 11; #1 b = 12;
		#1 b = 13; #1 b = 14; #1 b = 15;
		
		#1 a = 10; b = 0;
		#1 b = 1; #1 b = 2; #1 b = 3; #1 b = 4;
		#1 b = 5; #1 b = 6; #1 b = 7; #1 b = 8;
		#1 b = 9; #1 b = 10; #1 b = 11; #1 b = 12;
		#1 b = 13; #1 b = 14; #1 b = 15;
		
		#1 a = 11; b = 0;
		#1 b = 1; #1 b = 2; #1 b = 3; #1 b = 4;
		#1 b = 5; #1 b = 6; #1 b = 7; #1 b = 8;
		#1 b = 9; #1 b = 10; #1 b = 11; #1 b = 12;
		#1 b = 13; #1 b = 14; #1 b = 15;
		
		#1 a = 12; b = 0;
		#1 b = 1; #1 b = 2; #1 b = 3; #1 b = 4;
		#1 b = 5; #1 b = 6; #1 b = 7; #1 b = 8;
		#1 b = 9; #1 b = 10; #1 b = 11; #1 b = 12;
		#1 b = 13; #1 b = 14; #1 b = 15;
		
		#1 a = 13; b = 0;
		#1 b = 1; #1 b = 2; #1 b = 3; #1 b = 4;
		#1 b = 5; #1 b = 6; #1 b = 7; #1 b = 8;
		#1 b = 9; #1 b = 10; #1 b = 11; #1 b = 12;
		#1 b = 13; #1 b = 14; #1 b = 15;
		
		#1 a = 14; b = 0;
		#1 b = 1; #1 b = 2; #1 b = 3; #1 b = 4;
		#1 b = 5; #1 b = 6; #1 b = 7; #1 b = 8;
		#1 b = 9; #1 b = 10; #1 b = 11; #1 b = 12;
		#1 b = 13; #1 b = 14; #1 b = 15;
		
		#1 a = 15; b = 0;
		#1 b = 1; #1 b = 2; #1 b = 3; #1 b = 4;
		#1 b = 5; #1 b = 6; #1 b = 7; #1 b = 8;
		#1 b = 9; #1 b = 10; #1 b = 11; #1 b = 12;
		#1 b = 13; #1 b = 14; #1 b = 15;
	end
endmodule //principal