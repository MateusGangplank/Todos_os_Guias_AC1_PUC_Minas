// ---------------------
// guia02-Exercicio01
// Nome: Larissa Fernandes Leijoto
// Matricula: 410476
// ---------------------

// ---------------------
// -- NAND gate
// ---------------------

   module  Exercicio01(s4, a, b, c);
	output s4;
	input a, b, c;
	assign s4 = ~ (a & b & c);
	
   endmodule

   module testeMNAND;
	reg a, b, c;
	wire s1, s2, s3, s4;
                                          // SE POSSIVEL, DEFINIR EM OUTRO MODULO
	Exercicio01 MNAND1 (s1, a, a, a);
	Exercicio01 MNAND2 (s2, b, b, b);
	Exercicio01 MNAND3 (s3, c, c, c);
	Exercicio01 MNAND4 (s4, s1, s2, s3);

	initial begin
		a = 0;b = 0;c = 0;
	end

	initial begin

   #1 $display (" Larissa Fernandes Leijoto - 410476 ");
   #1 $display (" a | b | c = s4 ");
	
	$monitor (" %b | %b | %b = %b ", a,b,c,s4);
	   #1 a=0;b=0;c=1;
      #1 a=0;b=1;c=0;
      #1 a=0;b=1;c=1;
		#1 a=1;b=0;c=0;
		#1 a=1;b=0;c=1;
		#1 a=1;b=1;c=0;
		#1 a=1;b=1;c=1;
	end	
endmodule
