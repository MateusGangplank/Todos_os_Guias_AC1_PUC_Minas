// Nome: Felipe Torres
// Matricula: 412738

module andgate(output s, input a, input b, input c);
 assign s = (a & b) & c;
endmodule

module teste;
 reg x,y,w;
 wire z;
 
 andgate AND1 (z,x,y,w);
 
 initial begin
  x=0; y=0; w=0;
  $display("Teste\nx y w z");
  $monitor("%b %b %b %b",x,y,w,z);
  
  #1 x=0; y=0; w=1;
  #1 x=0; y=1; w=0;
  #1 x=0; y=1; w=1;
  #1 x=1; y=0; w=0;
  #1 x=1; y=0; w=1;
  #1 x=1; y=1; w=0;
  #1 x=1; y=1; w=1;
 end
 
endmodule