// Guia 05
// Nome: Raphaela Fernanda Silva
// Matricula: 420141


module operadorMD ( s0, s1, a, b);
output s0, s1;
input a, b;
wire s2;

xor XOR1(s0,a,b);
not NOT1(s2,a);
and AND1(s1,s2,b);

endmodule

module operadorDC ( s0, s1, a, b, v1 );
output s0, s1;
input a, b, v1;
wire s2, s3, s4;

operadorMD MD1(s2,s3,a,b);
operadorMD MD2(s4,s0,s2,v1);
or OR1(s1,s3,s4);

endmodule

module DC3Bits ( s, a, b);
output[3:0]s;
input[2:0]a,b;
wire[1:0]c;

operadorMD MD1(s[0],c[0],a[0],b[0]);
operadorDC DC1(s[1],c[1],a[1],b[1],c[0]);
operadorDC DC2(s[2],s[3],a[2],b[2],c[1]);

endmodule


module testDC;
reg[2:0]a,b;
wire[3:0]s;
integer i,j;

DC3Bits DC3B(s,a,b);

initial begin : start

a=0; b=0;

end

initial begin : main

#1 $display ( " Operador Diferen�a Completa - 3 Bits " );
#1 $display ( "   a  -  b   =  s   " );
	$monitor ( " %3b  %3b  = %4b ",a,b,s);
	
	for ( i = 0; i < 16; i = i + 1)begin
	 a = i;
	for ( j = 0; j < 16; j = j + 1)begin
	#1 b = j;
	end
	end
				
end

endmodule

/* Operador Diferen�a Completa - 3 Bits 
       a  -  b   =  s   
     000  000  = 0000 
     000  001  = 1111 
     000  010  = 1100 
     000  011  = 1101 
     000  100  = 1000 
     000  101  = 1011 
     000  110  = 1000 
     000  111  = 1001 
     000  000  = 0000 
     000  001  = 1111 
     000  010  = 1100 
     000  011  = 1101 
     000  100  = 1000 
     000  101  = 1011 
     000  110  = 1000 
     001  111  = 1000 
     001  000  = 0001 
     001  001  = 0000 
     001  010  = 1101 
     001  011  = 1100 
     001  100  = 1001 
     001  101  = 1000 
     001  110  = 1001 
     001  111  = 1000 
     001  000  = 0001 
     001  001  = 0000 
     001  010  = 1101 
     001  011  = 1100 
     001  100  = 1001 
     001  101  = 1000 
     001  110  = 1001 
     010  111  = 1011 
     010  000  = 1100 
     010  001  = 0001 
     010  010  = 0000 
     010  011  = 1111 
     010  100  = 1000 
     010  101  = 1001 
     010  110  = 1000 
     010  111  = 1011 
     010  000  = 1100 
     010  001  = 0001 
     010  010  = 0000 
     010  011  = 1111 
     010  100  = 1000 
     010  101  = 1001 
     010  110  = 1000 
     011  111  = 1000 
     011  000  = 1101 
     011  001  = 1100 
     011  010  = 0001 
     011  011  = 0000 
     011  100  = 1001 
     011  101  = 1000 
     011  110  = 1001 
     011  111  = 1000 
     011  000  = 1101 
     011  001  = 1100 
     011  010  = 0001 
     011  011  = 0000 
     011  100  = 1001 
     011  101  = 1000 
     011  110  = 1001 
     100  111  = 1101 
     100  000  = 1000 
     100  001  = 0011 
     100  010  = 0000 
     100  011  = 0001 
     100  100  = 0000 
     100  101  = 1111 
     100  110  = 1100 
     100  111  = 1101 
     100  000  = 1000 
     100  001  = 0011 
     100  010  = 0000 
     100  011  = 0001 
     100  100  = 0000 
     100  101  = 1111 
     100  110  = 1100 
     101  111  = 1100 
     101  000  = 1001 
     101  001  = 1000 
     101  010  = 0001 
     101  011  = 0000 
     101  100  = 0001 
     101  101  = 0000 
     101  110  = 1101 
     101  111  = 1100 
     101  000  = 1001 
     101  001  = 1000 
     101  010  = 0001 
     101  011  = 0000 
     101  100  = 0001 
     101  101  = 0000 
     101  110  = 1101 
     110  111  = 1111 
     110  000  = 0000 
     110  001  = 1001 
     110  010  = 1000 
     110  011  = 0011 
     110  100  = 1100 
     110  101  = 0001 
     110  110  = 0000 
     110  111  = 1111 
     110  000  = 0000 
     110  001  = 1001 
     110  010  = 1000 
     110  011  = 0011 
     110  100  = 1100 
     110  101  = 0001 
     110  110  = 0000 
     111  111  = 0000 
     111  000  = 0001 
     111  001  = 0000 
     111  010  = 1001 
     111  011  = 1000 
     111  100  = 1101 
     111  101  = 1100 
     111  110  = 0001 
     111  111  = 0000 
     111  000  = 0001 
     111  001  = 0000 
     111  010  = 1001 
     111  011  = 1000 
     111  100  = 1101 
     111  101  = 1100 
     111  110  = 0001 
     000  111  = 1001 
     000  000  = 0000 
     000  001  = 1111 
     000  010  = 1100 
     000  011  = 1101 
     000  100  = 1000 
     000  101  = 1011 
     000  110  = 1000 
     000  111  = 1001 
     000  000  = 0000 
     000  001  = 1111 
     000  010  = 1100 
     000  011  = 1101 
     000  100  = 1000 
     000  101  = 1011 
     000  110  = 1000 
     001  111  = 1000 
     001  000  = 0001 
     001  001  = 0000 
     001  010  = 1101 
     001  011  = 1100 
     001  100  = 1001 
     001  101  = 1000 
     001  110  = 1001 
     001  111  = 1000 
     001  000  = 0001 
     001  001  = 0000 
     001  010  = 1101 
     001  011  = 1100 
     001  100  = 1001 
     001  101  = 1000 
     001  110  = 1001 
     010  111  = 1011 
     010  000  = 1100 
     010  001  = 0001 
     010  010  = 0000 
     010  011  = 1111 
     010  100  = 1000 
     010  101  = 1001 
     010  110  = 1000 
     010  111  = 1011 
     010  000  = 1100 
     010  001  = 0001 
     010  010  = 0000 
     010  011  = 1111 
     010  100  = 1000 
     010  101  = 1001 
     010  110  = 1000 
     011  111  = 1000 
     011  000  = 1101 
     011  001  = 1100 
     011  010  = 0001 
     011  011  = 0000 
     011  100  = 1001 
     011  101  = 1000 
     011  110  = 1001 
     011  111  = 1000 
     011  000  = 1101 
     011  001  = 1100 
     011  010  = 0001 
     011  011  = 0000 
     011  100  = 1001 
     011  101  = 1000 
     011  110  = 1001 
     100  111  = 1101 
     100  000  = 1000 
     100  001  = 0011 
     100  010  = 0000 
     100  011  = 0001 
     100  100  = 0000 
     100  101  = 1111 
     100  110  = 1100 
     100  111  = 1101 
     100  000  = 1000 
     100  001  = 0011 
     100  010  = 0000 
     100  011  = 0001 
     100  100  = 0000 
     100  101  = 1111 
     100  110  = 1100 
     101  111  = 1100 
     101  000  = 1001 
     101  001  = 1000 
     101  010  = 0001 
     101  011  = 0000 
     101  100  = 0001 
     101  101  = 0000 
     101  110  = 1101 
     101  111  = 1100 
     101  000  = 1001 
     101  001  = 1000 
     101  010  = 0001 
     101  011  = 0000 
     101  100  = 0001 
     101  101  = 0000 
     101  110  = 1101 
     110  111  = 1111 
     110  000  = 0000 
     110  001  = 1001 
     110  010  = 1000 
     110  011  = 0011 
     110  100  = 1100 
     110  101  = 0001 
     110  110  = 0000 
     110  111  = 1111 
     110  000  = 0000 
     110  001  = 1001 
     110  010  = 1000 
     110  011  = 0011 
     110  100  = 1100 
     110  101  = 0001 
     110  110  = 0000 
     111  111  = 0000 
     111  000  = 0001 
     111  001  = 0000 
     111  010  = 1001 
     111  011  = 1000 
     111  100  = 1101 
     111  101  = 1100 
     111  110  = 0001 
     111  111  = 0000 
     111  000  = 0001 
     111  001  = 0000 
     111  010  = 1001 
     111  011  = 1000 
     111  100  = 1101 
     111  101  = 1100 
     111  110  = 0001 
     111  111  = 0000
*/



