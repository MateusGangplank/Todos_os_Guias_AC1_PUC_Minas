//-----
//Exercicio 05
//Andre Campolina
//381217
//-----

//-----
//porta nor de morgan
//-----

module norgate (output s, input p, input q);
	assign s=((~p)&(~q));
endmodule //norgate

//----
//tabela verdade
//----

module testnor;
	reg a, b;
	wire s;
	
	norgate NOR1(s, a, b);
	
	initial begin:start
		a=0; b=0;
	end
	
	initial begin
		$display("Exercicio05 - Andre Campolina - 381217");
		$display("Tabela Verdade porta NOR de morgan");
		$display("\na b\ts\n");
		$monitor("%b %b\t%b",a,b,s);
		#1 b=1;
		#1 a=1; b=0;
		#1 b=1;
	end
endmodule //testnor