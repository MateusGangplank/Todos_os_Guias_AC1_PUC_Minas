// Exercicio 001 � RAM 1X4
// Nome: �tila Martins Silva J�nior
// Matricula: 449014

module jkff(q,q1,j,k,c);
output q,q1;
input j,k,c;
reg q,q1;
initial begin q=1'b0; q1=1'b1; end
always @ (posedge c)
  begin
	case({j,k})
		 {1'b0,1'b0}:begin q=q; q1=q1; end
		 {1'b0,1'b1}: begin q=1'b0; q1=1'b1; end
		 {1'b1,1'b0}:begin q=1'b1; q1=1'b0; end
		 {1'b1,1'b1}: begin q=~q; q1=~q1; end
	endcase
   end
endmodule

module ram1x4(output[3:0] saida, input[3:0] ent, input clk, input rw, input addr);
	wire a1, a2, a3,s0, s1, s2, n0, n1, n2, n3, rw1;
	not(n0, ent[0]);
	not(n1, ent[1]);
	not(n2, ent[2]);
	not(n3, ent[3]);
	
	and(a1, clk, rw);
	and(a2, a1, addr);
	
	jkff JK0(s0,, ent[0], n0, a2);
	jkff JK1(s1,, ent[1], n1, a2);
	jkff JK2(s2,, ent[2], n2, a2);
	jkff JK3(s3,, ent[3], n3, a2);
	
	and(saida[0], addr, s0);
	and(saida[1], addr, s1);
	and(saida[2], addr, s2);
	and(saida[3], addr, s3);
endmodule

module testRam1x4;
	reg[3:0] entrada;
	reg clock, rw, addr;
	wire[3:0] saida;

	ram1x4 RAM1X4(saida, entrada, clock, rw, addr);
	
	initial begin
		$display("Exercicio01 - �tila Martins Silva J�nior - 449014");
		
		clock = 0; rw = 0; addr = 0; entrada = 4'b0000;
		
		$monitor("input: %b addr: %b rw: %b output: %b",entrada,addr,rw,saida);
		#4entrada = 4'b1111; 
		#4rw = 1; addr = 1; clock = 1;
		#4entrada = 4'b0101; 
		#4clock = 0;
		#4rw = 1; addr = 1; clock = 1;
		
		
		
	end
endmodule