// Nome: Caio Ragacci Pimentel
// Matr�cula: 405794

module metodoprovai ( saida,a,b,c,d );

output saida;
input a,b,c,d;
wire temp1,temp2,temp3,temp4,temp5,temp6,temp7,temp8,temp9,temp10;


xor XOR1 (temp1,a,d);
and AND1 (temp2,temp1,c);
xor XOR2 (temp3,a,b);
and AND2 (temp4,temp3,d);
not NOT1 (temp5,c);
and AND3 (temp6,b,temp5);
not NOT2 (temp7,d);
and AND4 (temp8,c,temp7);
or OR1   (temp9,temp6,temp8);
and AND5 (temp10,a,temp9);
or OR2   (saida,temp2,temp4,temp10);

endmodule
 
module testprova1;
reg a,b,c,d;
wire saida;

metodoprovai PROVAI ( saida,a,b,c,d );

initial begin:start
        a=0; b=0; c=0; d=0;
end

initial begin: main
#1 $display (" Circuito da questao i da prova ");
#1 $display (" a |  b |  c |  d  =  saida ");
  $monitor (" %b  | %b  | %b |  %b  =   %b ",a,b,c,d,saida);
           #1 a=0;    b=0;   c=0;   d=1;
			  #1 a=0;    b=0;   c=1;   d=0;
			  #1 a=0;    b=0;   c=1;   d=1;
			  #1 a=0;    b=1;   c=0;   d=0;
			  #1 a=0;    b=1;   c=0;   d=1;
			  #1 a=0;    b=1;   c=1;   d=0;
			  #1 a=0;    b=1;   c=1;   d=1;
			  #1 a=1;    b=0;   c=0;   d=0;
			  #1 a=1;    b=0;   c=0;   d=1;
			  #1 a=1;    b=0;   c=1;   d=0;
			  #1 a=1;    b=0;   c=1;   d=1;
			  #1 a=1;    b=1;   c=0;   d=0;
			  #1 a=1;    b=1;   c=0;   d=1;
			  #1 a=1;    b=1;   c=1;   d=0;
			  #1 a=1;    b=1;   c=1;   d=1;
			  
			  
			  
end
endmodule
