// ------------------------- 
// Exemplo0041 - FULL ADDER 
// Nome:Mateus Guilherme do Carmo Cruz
// Matricula: 427446
// ------------------------- 
 `include "FullAdder.v"

module test_fullAdder; 
// ------------------------- definir dados 
	reg [3:0] x; 
	reg [3:0] y; 
	reg carry; 
	wire [3:0] soma;
	
// ------------------------- inst�ncia
	fullAdder4bits fa1(soma,x,y, 0);
	
// ------------------------- parte principal 
	initial begin 
		$display("Exemplo0041 - Mateus Guilherme do Carmo Cruz - 427446"); 
		$display("Test ALU's full adder"); 
		x = 4'b0000;
		y = 4'b0000;
		carry = 0;
		$display("\t  \tt\tx + y = soma");
		$monitor("%d %4b + %4b = %4b",$time,x,y,soma);
		#1 y = 4'b0001;
		#1 y = 4'b0010;
		#1 y = 4'b0011;
		#1 y = 4'b0100;
		#1 y = 4'b0101;
		#1 y = 4'b0110;
		#1 y = 4'b0111;
		#1 y = 4'b1000;
		#1 y = 4'b1001;
		#1 y = 4'b1010;
		#1 y = 4'b1011;
		#1 y = 4'b1100;
		#1 y = 4'b1101;
		#1 y = 4'b1110;
		#1 y = 4'b1111;
		
		#1 x = 4'b0001; y = 4'b0000;
		#1 y = 4'b0001;
		#1 y = 4'b0010;
		#1 y = 4'b0011;
		#1 y = 4'b0100;
		#1 y = 4'b0101;
		#1 y = 4'b0110;
		#1 y = 4'b0111;
		#1 y = 4'b1000;
		#1 y = 4'b1001;
		#1 y = 4'b1010;
		#1 y = 4'b1011;
		#1 y = 4'b1100;
		#1 y = 4'b1101;
		#1 y = 4'b1110;
		#1 y = 4'b1111;
		
		#1 x = 4'b0010; y = 4'b0000;
		#1 y = 4'b0001;
		#1 y = 4'b0010;
		#1 y = 4'b0011;
		#1 y = 4'b0100;
		#1 y = 4'b0101;
		#1 y = 4'b0110;
		#1 y = 4'b0111;
		#1 y = 4'b1000;
		#1 y = 4'b1001;
		#1 y = 4'b1010;
		#1 y = 4'b1011;
		#1 y = 4'b1100;
		#1 y = 4'b1101;
		#1 y = 4'b1110;
		#1 y = 4'b1111;
		
		#1 x = 4'b1000; y = 4'b0000;
		#1 y = 4'b0001;
		#1 y = 4'b0010;
		#1 y = 4'b0011;
		#1 y = 4'b0100;
		#1 y = 4'b0101;
		#1 y = 4'b0110;
		#1 y = 4'b0111;
		#1 y = 4'b1000;
		#1 y = 4'b1001;
		#1 y = 4'b1010;
		#1 y = 4'b1011;
		#1 y = 4'b1100;
		#1 y = 4'b1101;
		#1 y = 4'b1110;
		#1 y = 4'b1111;
		
		#1 x = 4'b1101; y = 4'b0000;
		#1 y = 4'b0001;
		#1 y = 4'b0010;
		#1 y = 4'b0011;
		#1 y = 4'b0100;
		#1 y = 4'b0101;
		#1 y = 4'b0110;
		#1 y = 4'b0111;
		#1 y = 4'b1000;
		#1 y = 4'b1001;
		#1 y = 4'b1010;
		#1 y = 4'b1011;
		#1 y = 4'b1100;
		#1 y = 4'b1101;
		#1 y = 4'b1110;
		#1 y = 4'b1111;
		
		#1 x = 4'b1111; y = 4'b0000;
		#1 y = 4'b0001;
		#1 y = 4'b0010;
		#1 y = 4'b0011;
		#1 y = 4'b0100;
		#1 y = 4'b0101;
		#1 y = 4'b0110;
		#1 y = 4'b0111;
		#1 y = 4'b1000;
		#1 y = 4'b1001;
		#1 y = 4'b1010;
		#1 y = 4'b1011;
		#1 y = 4'b1100;
		#1 y = 4'b1101;
		#1 y = 4'b1110;
		#1 y = 4'b1111;
	end 
endmodule // test_fullAdder 