// ---------------------
// Guia05
// Nome: Lucas Teixeira Santos
// Matricula: 415383
// ---------------------

// ---------------------
// -- test ex01
// -- Expressao Simplificada:
// -- S = a ^ b
// -- C = a & b
// ---------------------

module meiasoma (a,b,s0,s1);
 output s0,s1;
 input  a, b;
 assign s1 = a & b;
 xor XOR (s0,a,b);
         
endmodule  // fim modulo principal

module somacompleta(a,b,cin,s0,s1);
output s0,s1;
input a,b,cin;
wire c1,c2;
meiasoma HA (cin,a,s,c1);
meiasoma HA2 (s,b,s0,c2);
assign s1 = c1 | c2;
endmodule
    
module testex1;
reg [2:0]a;
reg [2:0]b;
wire c0,s0,s1,c1,s2,c2;
meiasoma HA (a[0],b[0],s0,c0);
somacompleta FA (a[1],b[1],c0,s1,c1);
somacompleta FA2 (a[2],b[2],c1,s2,c2);
initial begin
      $display("Exercicio 01 - Lucas Teixeira Santos - 415383");
      $display("Soma Completa 3 Bits.");
      $display("AAA  +  BBB  =  CCCC");
a = 3'b000;
b = 3'b000;
   #1	 $monitor("%b  +  %b  =  %b%b%b%b", a, b, c2,s2,s1,s0);
   #1  b=b+1;
   #1  b=b+1;
	#1  b=b+1;
	#1  b=b+1;
   #1  b=b+1;
   #1  b=b+1;
	#1  b=b+1;
	#1  a=a+1; b=0;
	#1  b=b+1;
   #1  b=b+1;
   #1  b=b+1;
	#1  b=b+1;
	#1  b=b+1;
   #1  b=b+1;
   #1  b=b+1;
	#1  a=a+1; b=0;	
	#1  b=b+1;
   #1  b=b+1;
   #1  b=b+1;
	#1  b=b+1;
	#1  b=b+1;
   #1  b=b+1;
   #1  b=b+1;
	#1  a=a+1; b=0;
	#1  b=b+1;
   #1  b=b+1;
   #1  b=b+1;
	#1  b=b+1;
	#1  b=b+1;
   #1  b=b+1;
   #1  b=b+1;
	#1  a=a+1; b=0;
	#1  b=b+1;
   #1  b=b+1;
   #1  b=b+1;
	#1  b=b+1;
	#1  b=b+1;
   #1  b=b+1;
   #1  b=b+1;
	#1  a=a+1; b=0;
	#1  b=b+1;
   #1  b=b+1;
   #1  b=b+1;
	#1  b=b+1;
	#1  b=b+1;
   #1  b=b+1;
   #1  b=b+1;
	#1  a=a+1; b=0;	
	#1  b=b+1;
   #1  b=b+1;
   #1  b=b+1;
	#1  b=b+1;
	#1  b=b+1;
   #1  b=b+1;
   #1  b=b+1;
	#1  a=a+1; b=0;	
	#1  b=b+1;
   #1  b=b+1;
   #1  b=b+1;
	#1  b=b+1;
	#1  b=b+1;
   #1  b=b+1;
   #1  b=b+1;
 end

endmodule 
/* test
    Soma Completa 3 Bits.
    AAA  +  BBB  =  CCCC
    000  +  000  =  0000
    000  +  001  =  0001
    000  +  010  =  0010
    000  +  011  =  0011
    000  +  100  =  0100
    000  +  101  =  0101
    000  +  110  =  0110
    000  +  111  =  0111
    001  +  000  =  0001
    001  +  001  =  0010
    001  +  010  =  0011
    001  +  011  =  0100
    001  +  100  =  0101
    001  +  101  =  0110
    001  +  110  =  0111
    001  +  111  =  1000
    010  +  000  =  0010
    010  +  001  =  0011
    010  +  010  =  0100
    010  +  011  =  0101
    010  +  100  =  0110
    010  +  101  =  0111
    010  +  110  =  1000
    010  +  111  =  1001
    011  +  000  =  0011
    011  +  001  =  0100
    011  +  010  =  0101
    011  +  011  =  0110
    011  +  100  =  0111
    011  +  101  =  1000
    011  +  110  =  1001
    011  +  111  =  1010
    100  +  000  =  0100
    100  +  001  =  0101
    100  +  010  =  0110
    100  +  011  =  0111
    100  +  100  =  1000
    100  +  101  =  1001
    100  +  110  =  1010
    100  +  111  =  1011
    101  +  000  =  0101
    101  +  001  =  0110
    101  +  010  =  0111
    101  +  011  =  1000
    101  +  100  =  1001
    101  +  101  =  1010
    101  +  110  =  1011
    101  +  111  =  1100
    110  +  000  =  0110
    110  +  001  =  0111
    110  +  010  =  1000
    110  +  011  =  1001
    110  +  100  =  1010
    110  +  101  =  1011
    110  +  110  =  1100
    110  +  111  =  1101
    111  +  000  =  0111
    111  +  001  =  1000
    111  +  010  =  1001
    111  +  011  =  1010
    111  +  100  =  1011
    111  +  101  =  1100
    111  +  110  =  1101
    111  +  111  =  1110
/*