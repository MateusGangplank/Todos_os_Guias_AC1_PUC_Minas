// ---------------------
// PUC-Minas - Instituto de Inform�tica
// ARQ1 Guia-03 Exercicio 03
// Data de entrega: 14-18/02/2011
// Nome: Pedro Tronbin
// Matricula: 410473
// ---------------------


// ---------------------
// -- test ex 03
// ---------------------

 module testex03;
 reg   a, b;
 wire  nOut, cOut, s, s0, s1, s2, nand4, nand5, notA, notB, snotAANDb, saANDnotB, notC;
 
 nand NAND2 (notA, a, a); // ~A.
 nand NAND3 (notB, b, b); // ~B.
 nand NAND4 (saANDnotB, a, notB); // (A&~B)
 nand NAND5 (snotAANDb, notA, b);  //(~A&B)
 nand NAND6 (nand4, saANDnotB, saANDnotB);  // ~
 nand NAND7 (nand5, snotAANDb, snotAANDb);  // ~
 nand NAND8 (s2, nand4, nand5);      
 nand NAND9 (s1, nand4, s2);         
 nand NAND10(s0, nand5, s2);        
 nand NAND11(s, s0, s1);            
 nand NAND0 (nOut, notC, b);  // no carry out
 nand NANDX (notC, a, a);
 nand NAND1 (cOut, nOut, nOut);  // carry out
          
         
 initial begin
 
      $display("Exercicio 03 - Pedro Tronbin - 410473");
      $display("Half Subtractor Test.");
      $display("A  -  B  =  C  S");
		
      a=0; b=0;
		 
  	#1	 $monitor("%b  -  %b  =  %b  %b", a, b, cOut, s);
   #1  a=0; b=1;
   #1  a=1; b=0;
   #1  a=1; b=1;
 
 end

endmodule // testex03

/* SAIDA

Exercicio 03 - Pedro Tronbin - 410473
    Half Subtractor Test.
    A  -  B  =  C  S
    0  -  0  =  0  0
    0  -  1  =  1  1
    1  -  0  =  0  1
    1  -  1  =  0  0

