// --------------------- 
// Exercicio01-05 - NOR
// Nome: Lucas Siqueira Chagas	 
// Matricula: 380783
// --------------------- 
// --------------------- 
// -- NAND
// --------------------- 
module norgate (output s, 
input p, 
input q); 
assign s = ~p&~q; 
endmodule // norgate 
// --------------------- 
// -- test norgate 
// --------------------- 
module testnorgate; 
// ------------------------- dados locais 
reg a,b; // definir registrador 
wire s; // definir conexao (fio) 
// ------------------------- instancia 
norgate NOR1 (s, a, b); 
// ------------------------- preparacao 
initial begin:start 
a=0; 
b=0;
end 
// ------------------------- parte principal 
initial begin:main 
$display("Exercicio01-05 - Lucas Siqueira Chagas - 380783"); 
$display("Test NOR gate por de morgan"); 
$display("\n (~a & ~b) = s\n"); 
a=0; b=0;
$monitor("(~%b & ~%b) = %b", a, b, s);
#1 a=0; b=1;
#1 a=1; b=0;
#1 a=1; b=1;
end 
endmodule // testnorgate 