// -------------------------
// Exemplo0018 - Exercicio03 
// Nome: Lorena Danielle Gon�alves Bento 
// Matricula: 435049
// ------------------------- 
// ------------------------- 
// test number system 
// ------------------------- 
// -- modulo --
module testexer03; 
// ------------------------- definir dados 
reg [4:0] a; 
reg [4:0] b; 
reg [9:0] c; 
reg [2:0] d; 
reg [3:0] e;
// ------------------------- parte principal 
initial begin:start
$display("Exercicio03 - Lorena Danielle Gon�alves Bento - 435049"); 
$display("Test number system"); 
a = ~6'o54 + 1;
b = ~5'h1B+1;
c = ~13 + 1;
d = ~5'h1B + 1;
e = 5'd25 + 1;
$display("\nResultado em binario");
$display("a = %d = %5b", a, a); 
$display("b = %d = %5b", b, b); 
$display("c = %d = %4b", c, c);
$display("d = %d = %4b", d, d);
$display("e = %d = %4b", e, e);
end 
endmodule // testexer03