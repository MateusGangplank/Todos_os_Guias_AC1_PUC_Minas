//
// Nome: Thaise Souto Martins
//

module Exer1 (s, s1, a, b);
input a, b;
output s, s1;

 xor XOR1 (s,a,b);
 and AND1 (s1,a,b);
 
endmodule 



module soma1 (s2, s4, a, b, c);
input a, b, c;
output  s2, s4;
wire s, s1, s3;

Exer1 Meia1 (s, s1, a, b);
Exer1 Meia2 (s2, s3, s, c);
or ou (s4, s1, s3);

endmodule  



module teste;
 reg   a, b, c, d, e ,f;
 wire  s, s1, s2, s3, s4, s5;
          
			 
			 
 Exer1 Meia3 (s,s1,c,f);
 soma1 Soma2 (s2, s3, s1, b, e);
 soma1 Soma3 (s4, s5, s3, a, d);



         
 initial begin
     	$display("Igor Rodrigues de Oliveira - 380771");
      $display("Exercicio 01");
		$display("AC - 2010");
      $display("\na b c  d e f   s");
 	   $monitor("%b %b %b  %b %b %b  %b%b%b | %b", a, b, c, d, e, f, s4, s2, s, s5);
 		
         a=0; b=0; c=0; d=0; e=0; f=0;
      #1 a=0; b=0; c=0; d=0; e=0; f=1;
		#1 a=0; b=0; c=0; d=0; e=1; f=0;
		#1 a=0; b=0; c=0; d=0; e=1; f=1;
		#1 a=0; b=0; c=0; d=1; e=0; f=0;
		#1 a=0; b=0; c=0; d=1; e=0; f=1;
		#1 a=0; b=0; c=0; d=1; e=1; f=0;
		#1 a=0; b=0; c=0; d=1; e=1; f=1;
		#1 a=0; b=0; c=1; d=0; e=0; f=0;
		#1 a=0; b=0; c=1; d=0; e=0; f=1;
		#1 a=0; b=0; c=1; d=0; e=1; f=0;
		#1 a=0; b=0; c=1; d=0; e=1; f=1;
		#1 a=0; b=0; c=1; d=1; e=0; f=0;
		#1 a=0; b=0; c=1; d=1; e=0; f=1;
		#1 a=0; b=0; c=1; d=1; e=1; f=0;
		#1 a=0; b=0; c=1; d=1; e=1; f=1;
		#1 a=0; b=1; c=0; d=0; e=0; f=0;
		#1 a=0; b=1; c=0; d=0; e=0; f=1;
		#1 a=0; b=1; c=0; d=0; e=1; f=0;
		#1 a=0; b=1; c=0; d=0; e=1; f=1;
		#1 a=0; b=1; c=0; d=1; e=0; f=0;
		#1 a=0; b=1; c=0; d=1; e=0; f=1;
		#1 a=0; b=1; c=0; d=1; e=1; f=0;
		#1 a=0; b=1; c=0; d=1; e=1; f=1;
		#1 a=0; b=1; c=1; d=0; e=0; f=0;
		#1 a=0; b=1; c=1; d=0; e=0; f=1;
		#1 a=0; b=1; c=1; d=0; e=1; f=0;
		#1 a=0; b=1; c=1; d=0; e=1; f=1;
		#1 a=0; b=1; c=1; d=1; e=0; f=0;
		#1 a=0; b=1; c=1; d=1; e=0; f=1;
		#1 a=0; b=1; c=1; d=1; e=1; f=0;
		#1 a=0; b=1; c=1; d=1; e=1; f=1;
		#1 a=1; b=1; c=0; d=0; e=0; f=0;
		#1 a=1; b=0; c=0; d=0; e=0; f=1;
		#1 a=1; b=0; c=0; d=0; e=1; f=0;
		#1 a=1; b=0; c=0; d=0; e=1; f=1;
		#1 a=1; b=0; c=0; d=1; e=0; f=0;
		#1 a=1; b=0; c=0; d=1; e=0; f=1;
		#1 a=1; b=0; c=0; d=1; e=1; f=0;
		#1 a=1; b=0; c=0; d=1; e=1; f=1;
		#1 a=1; b=0; c=1; d=0; e=0; f=0;
		#1 a=1; b=0; c=1; d=0; e=0; f=1;
		#1 a=1; b=0; c=1; d=0; e=1; f=0;
		#1 a=1; b=0; c=1; d=0; e=1; f=1;
		#1 a=1; b=0; c=1; d=1; e=0; f=0;
		#1 a=1; b=0; c=1; d=1; e=0; f=1;
		#1 a=1; b=0; c=1; d=1; e=1; f=0;
		#1 a=1; b=0; c=1; d=1; e=1; f=1;
		#1 a=1; b=1; c=0; d=0; e=0; f=0;
		#1 a=1; b=1; c=0; d=0; e=0; f=1;
		#1 a=1; b=1; c=0; d=0; e=1; f=0;
		#1 a=1; b=1; c=0; d=0; e=1; f=1;
		#1 a=1; b=1; c=0; d=1; e=0; f=0;
		#1 a=1; b=1; c=0; d=1; e=0; f=1;
		#1 a=1; b=1; c=0; d=1; e=1; f=0;
		#1 a=1; b=1; c=0; d=1; e=1; f=1;
		#1 a=1; b=1; c=1; d=0; e=0; f=0;
		#1 a=1; b=1; c=1; d=0; e=0; f=1;
		#1 a=1; b=1; c=1; d=0; e=1; f=0;
		#1 a=1; b=1; c=1; d=0; e=1; f=1;
		#1 a=1; b=1; c=1; d=1; e=0; f=0;
		#1 a=1; b=1; c=1; d=1; e=0; f=1;
		#1 a=1; b=1; c=1; d=1; e=1; f=0;
		#1 a=1; b=1; c=1; d=1; e=1; f=1;
		
 end

endmodule