// -------------------------
// Exemplo0034 - F4
// Nome: Davidson Francis
// Matricula: 466499
// -------------------------


// -------------------------
// f4_gate
// -------------------------

module f4 (output s,
           input  a,
           input  b,
           input  c1, input c2);

wire temp[0:8];

 or   OR1  (temp[0], a,b);
 nor  NOR1 (temp[1], a,b);
 xor  XOR1 (temp[2], a,b);
 xnor XNOR1(temp[3], a,b);
// USAR PORTA not PARA ~c1, ~c2 TAMBEM
 and AND1(temp[4],  ~c1,~c2,temp[0]);
 and AND2(temp[5],  ~c1, c2,temp[1]);
 and AND3(temp[6],   c1, c2,temp[2]);
 and AND4(temp[7],   c1, c2,temp[3]);

 or OR2(temp[8], temp[4],temp[5],temp[6],temp[7]);

 assign s = temp[8];

endmodule


module test_f4;

// ------------------------- definir dados
reg  a;
reg  b;
reg  c1;
reg  c2;
wire s;

f4 modulo (s, a,b,c1,c2);


initial begin:start
  a=0;b=0;  c1=0;c2=0;
end


// ------------------------- parte principal
initial begin:main
  $display("Exemplo0034 - Davidson Francis - 466499");
  $display("Test LU's module");
  
  $display("a  b  chave  saida");
  $monitor("%b  %b  %b %b     %b", a,b,c1,c2, s);
 
  #1 a = 0; b = 0;   c1 = 0; c2=0;
  #1 a = 0; b = 0;   c1 = 0; c2=1;
  #1 a = 0; b = 0;   c1 = 1; c2=0;
  #1 a = 0; b = 0;   c1 = 1; c2=1;
  #1 a = 0; b = 1;   c1 = 0; c2=0;
  #1 a = 0; b = 1;   c1 = 0; c2=1;
  #1 a = 0; b = 1;   c1 = 1; c2=0;
  #1 a = 0; b = 1;   c1 = 1; c2=1;
  
  #1 a = 1; b = 0;   c1 = 0; c2=0;
  #1 a = 1; b = 0;   c1 = 0; c2=1;
  #1 a = 1; b = 0;   c1 = 1; c2=0;
  #1 a = 1; b = 0;   c1 = 1; c2=1;
  #1 a = 1; b = 1;   c1 = 0; c2=0;
  #1 a = 1; b = 1;   c1 = 0; c2=1;
  #1 a = 1; b = 1;   c1 = 1; c2=0;
  #1 a = 1; b = 1;   c1 = 1; c2=1;
end
endmodule
