// ---------------------------
// -- CLOCK Generator
// Herbert Alves Batista - 461971
// ---------------------------
module clock ( clk );
output clk;
reg clk;
initial
begin
clk = 1'b0;
end
always
begin
#12 clk = ~clk;
end
endmodule // clock ( )
module Exemplo0044;
wire clk;
clock CLK1 ( clk );
initial begin
$dumpfile ( "Exemplo0041.vcd" );
$dumpvars;
#120 $finish;
end
endmodule // Exemplo044 ( )