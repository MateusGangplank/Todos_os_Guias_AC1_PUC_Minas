// ------------------------- 
// Exemplo0004 - OR 
// Nome: Gabriel Luiz M. G. Vieira 
// Matricula: 441691 
// ------------------------- 
// ------------------------- 
// -- or gate 
// ------------------------- 
module orgate ( output s, 
input p, q); 
assign s = p | q; 
endmodule // orgate 
// --------------------- 
// -- test or gate 
// --------------------- 
module testorgate; 
// ------------------------- dados locais 
reg a, b; // definir registradores 
wire s; // definir conexao (fio) 
// ------------------------- instancia 
orgate OR1 (s, a, b); 
// ------------------------- preparacao 
initial begin:start 
// atribuicao simultanea 
// dos valores iniciais 
a=0; b=0; 
end 
// ------------------------- parte principal 
initial begin 
$display("Exemplo0004 - Gabriel Luiz M. G. Vieira - 441691"); 
$display("Test OR gate"); 
$display("\na | b = s\n"); 
$monitor("%b & %b = %b", a, b, s); 
#1a=0; b=0;  
#1a=0; b=1; 
#1a=1; b=0; 
#1a=1; b=1; 
end 
endmodule // testorgate 