//ARQ1 - Guia07 - Eduardo Botelho de Andrade

`include "mealy.v"
`include "moore.v"

module ex0701;
 reg clk,reset,x;
 wire m1,m2;
 
 mealy mealy1 (m1,x,clk,reset);
 moore moore1 (m2,x,clk,reset);
 
 initial
  begin
   $display("Time    X     Mealy  Moore");
   
   //initial values
    clk = 1;
    reset = 0;
    x = 0;
   
  //input signal changing
  

  // input signal changing
    #5    reset = 1; 
    #10  x = 1; 
    #10  x = 0; 
    #10  x = 1; 
    #20  x = 0; 
    #10  x = 1; 
    #10  x = 1; 
    #10  x = 0;
    #10  x = 1;
 
    #30 $finish;
  end // initial

 always
  #5 clk = ~clk;

 always @( posedge clk ) 
  begin 
   $display ("%4d  %4b  %4b %5b", $time, x, m1, m2);
  end // always at positive edge clocking changing
endmodule