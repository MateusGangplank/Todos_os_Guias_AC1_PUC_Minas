//ARQ1 - Eduardo Botelho de Andrade - Guia03
// -------------------------
// Exemplo0031 - F4


// Nome: xxx yyy zzz
// Matricula: 999999 
// ------------------------- 
 
// ------------------------- 
//  f4_gate 
// -------------------------
module f4 (output [3:0] s, 
           input  [3:0] a,
           input  [3:0] b); 
 
 and and1 (s[0],a[0],b[0]);
 and and2 (s[1],a[1],b[1]);
 and and3 (s[2],a[2],b[2]);
 and and4 (s[3],a[3],b[3]);
 
endmodule // f4 
 
module test_f4; 
// ------------------------- definir dados 
       reg  [3:0] x; 
       reg  [3:0] y; 
       wire [3:0] z; 
 
       f4 modulo (z, x, y); 
 
// ------------------------- parte principal 
 
   initial begin 
      $display("Eduardo Botelho de Andrade - 427395");
      $display("Test LU's module");
      $monitor("x = %b , y = %b , z = %b",x,y,z);

      #1 x = 4'b0000; y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;
      
      #1 x = 4'b0001;
      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;
      
      #1 x = 4'b0010;
      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;
      
      #1 x = 4'b0011;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;
      
      #1 x = 4'b0100;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;
      
      #1 x = 4'b0101;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;
      
      #1 x = 4'b0110;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;
      
      #1 x = 4'b0111;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;
      
      #1 x = 4'b1000; 

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;
      
      #1 x = 4'b1001;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;
      
      #1 x = 4'b1010;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;
      
      #1 x = 4'b1011;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;
      
      #1 x = 4'b1100;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;

      #1 x=4'b1101;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;

      #1 x=4'b1110;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;

      #1 x=4'b1111;

      #1 y = 4'b0000;
      #1 y = 4'b0001;
      #1 y = 4'b0010;
      #1 y = 4'b0011;
      #1 y = 4'b0100;
      #1 y = 4'b0101;
      #1 y = 4'b0110;
      #1 y = 4'b0111;
      #1 y = 4'b1000;
      #1 y = 4'b1001;
      #1 y = 4'b1010;
      #1 y = 4'b1011;
      #1 y = 4'b1100;
      #1 y = 4'b1101;
      #1 y = 4'b1111;

   end 
 
endmodule // test_f4 
